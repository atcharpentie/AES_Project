
module AES_top ( data_in, key_in, out_data, ready, rst, clk );
  input [127:0] data_in;
  input [127:0] key_in;
  output [127:0] out_data;
  input rst, clk;
  output ready;
  wire   n2995, n2996, n3125, n3126, n3127, n3128, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, U99_DATA1_0, U99_DATA1_1, U99_DATA1_2, U99_DATA1_3,
         U99_DATA1_4, U99_DATA1_5, U99_DATA1_6, U99_DATA1_7, U99_DATA1_8,
         U99_DATA1_9, U99_DATA1_10, U99_DATA1_11, U99_DATA1_12, U99_DATA1_13,
         U99_DATA1_14, U99_DATA1_15, U99_DATA1_16, U99_DATA1_17, U99_DATA1_18,
         U99_DATA1_19, U99_DATA1_20, U99_DATA1_21, U99_DATA1_22, U99_DATA1_23,
         U99_DATA1_24, U99_DATA1_25, U99_DATA1_26, U99_DATA1_27, U99_DATA1_28,
         U99_DATA1_29, U99_DATA1_30, U99_DATA1_31, U99_DATA1_32, U99_DATA1_33,
         U99_DATA1_34, U99_DATA1_35, U99_DATA1_36, U99_DATA1_37, U99_DATA1_38,
         U99_DATA1_39, U99_DATA1_40, U99_DATA1_41, U99_DATA1_42, U99_DATA1_43,
         U99_DATA1_44, U99_DATA1_45, U99_DATA1_46, U99_DATA1_47, U99_DATA1_48,
         U99_DATA1_49, U99_DATA1_50, U99_DATA1_51, U99_DATA1_52, U99_DATA1_53,
         U99_DATA1_54, U99_DATA1_55, U99_DATA1_56, U99_DATA1_57, U99_DATA1_58,
         U99_DATA1_59, U99_DATA1_60, U99_DATA1_61, U99_DATA1_62, U99_DATA1_63,
         U99_DATA1_64, U99_DATA1_65, U99_DATA1_66, U99_DATA1_67, U99_DATA1_68,
         U99_DATA1_69, U99_DATA1_70, U99_DATA1_71, U99_DATA1_72, U99_DATA1_73,
         U99_DATA1_74, U99_DATA1_75, U99_DATA1_76, U99_DATA1_77, U99_DATA1_78,
         U99_DATA1_79, U99_DATA1_80, U99_DATA1_81, U99_DATA1_82, U99_DATA1_83,
         U99_DATA1_84, U99_DATA1_85, U99_DATA1_86, U99_DATA1_87, U99_DATA1_88,
         U99_DATA1_89, U99_DATA1_90, U99_DATA1_91, U99_DATA1_92, U99_DATA1_93,
         U99_DATA1_94, U99_DATA1_95, U99_DATA1_96, U99_DATA1_97, U99_DATA1_98,
         U99_DATA1_99, U99_DATA1_100, U99_DATA1_101, U99_DATA1_102,
         U99_DATA1_103, U99_DATA1_104, U99_DATA1_105, U99_DATA1_106,
         U99_DATA1_107, U99_DATA1_108, U99_DATA1_109, U99_DATA1_110,
         U99_DATA1_111, U99_DATA1_112, U99_DATA1_113, U99_DATA1_114,
         U99_DATA1_115, U99_DATA1_116, U99_DATA1_117, U99_DATA1_118,
         U99_DATA1_119, U99_DATA1_120, U99_DATA1_121, U99_DATA1_122,
         U99_DATA1_123, U99_DATA1_124, U99_DATA1_125, U99_DATA1_126,
         U99_DATA1_127, U51_Z_0, U51_Z_1, U51_Z_2, U51_Z_3, U49_Z_0, U49_Z_1,
         U49_Z_2, U49_Z_3, U49_Z_4, U49_Z_5, U49_Z_6, U49_Z_7, U49_Z_8,
         U49_Z_9, U49_Z_10, U49_Z_11, U49_Z_12, U49_Z_13, U49_Z_14, U49_Z_15,
         U49_Z_16, U49_Z_17, U49_Z_18, U49_Z_19, U49_Z_20, U49_Z_21, U49_Z_22,
         U49_Z_23, U49_Z_24, U49_Z_25, U49_Z_26, U49_Z_27, U49_Z_28, U49_Z_29,
         U49_Z_30, U49_Z_31, U49_Z_32, U49_Z_33, U49_Z_34, U49_Z_35, U49_Z_36,
         U49_Z_37, U49_Z_38, U49_Z_39, U49_Z_40, U49_Z_41, U49_Z_42, U49_Z_43,
         U49_Z_44, U49_Z_45, U49_Z_46, U49_Z_47, U49_Z_48, U49_Z_49, U49_Z_50,
         U49_Z_51, U49_Z_52, U49_Z_53, U49_Z_54, U49_Z_55, U49_Z_56, U49_Z_57,
         U49_Z_58, U49_Z_59, U49_Z_60, U49_Z_61, U49_Z_62, U49_Z_63, U49_Z_64,
         U49_Z_65, U49_Z_66, U49_Z_67, U49_Z_68, U49_Z_69, U49_Z_70, U49_Z_71,
         U49_Z_72, U49_Z_73, U49_Z_74, U49_Z_75, U49_Z_76, U49_Z_77, U49_Z_78,
         U49_Z_79, U49_Z_80, U49_Z_81, U49_Z_82, U49_Z_83, U49_Z_84, U49_Z_85,
         U49_Z_86, U49_Z_87, U49_Z_88, U49_Z_89, U49_Z_90, U49_Z_91, U49_Z_92,
         U49_Z_93, U49_Z_94, U49_Z_95, U49_Z_96, U49_Z_97, U49_Z_98, U49_Z_99,
         U49_Z_100, U49_Z_101, U49_Z_102, U49_Z_103, U49_Z_104, U49_Z_105,
         U49_Z_106, U49_Z_107, U49_Z_108, U49_Z_109, U49_Z_110, U49_Z_111,
         U49_Z_112, U49_Z_113, U49_Z_114, U49_Z_115, U49_Z_116, U49_Z_117,
         U49_Z_118, U49_Z_119, U49_Z_120, U49_Z_121, U49_Z_122, U49_Z_123,
         U49_Z_124, U49_Z_125, U49_Z_126, U49_Z_127, U47_Z_1, U46_Z_1,
         r424_A_0_, r424_A_1_, r424_A_2_, r424_A_3_, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         R2_n2407, R2_n2406, R2_n2405, R2_n2404, R2_n2403, R2_n2402, R2_n2401,
         R2_n2400, R2_n2399, R2_n2398, R2_n2397, R2_n2396, R2_n2395, R2_n2394,
         R2_n2393, R2_n2392, R2_n2391, R2_n2390, R2_n2389, R2_n2388, R2_n2387,
         R2_n2386, R2_n2385, R2_n2384, R2_n2383, R2_n2382, R2_n2381, R2_n2380,
         R2_n2379, R2_n2378, R2_n2377, R2_n2376, R2_n2375, R2_n2374, R2_n2373,
         R2_n2372, R2_n2371, R2_n2370, R2_n2369, R2_n2368, R2_n2367, R2_n2366,
         R2_n2365, R2_n2364, R2_n2363, R2_n2362, R2_n2361, R2_n2360, R2_n2359,
         R2_n2358, R2_n2357, R2_n2356, R2_n2355, R2_n2354, R2_n2353, R2_n2352,
         R2_n2351, R2_n2350, R2_n2349, R2_n2348, R2_n2347, R2_n2346, R2_n2345,
         R2_n2344, R2_n2343, R2_n2342, R2_n2341, R2_n2340, R2_n2339, R2_n2338,
         R2_n2337, R2_n2336, R2_n2335, R2_n2334, R2_n2333, R2_n2332, R2_n2331,
         R2_n2330, R2_n2329, R2_n2328, R2_n2327, R2_n2326, R2_n2325, R2_n2324,
         R2_n2323, R2_n2322, R2_n2321, R2_n2320, R2_n2319, R2_n2318, R2_n2317,
         R2_n2316, R2_n2315, R2_n2314, R2_n2313, R2_n2312, R2_n2311, R2_n2310,
         R2_n2309, R2_n2308, R2_n2307, R2_n2306, R2_n2305, R2_n2304, R2_n2303,
         R2_n2302, R2_n2301, R2_n2300, R2_n2299, R2_n2298, R2_n2297, R2_n2296,
         R2_n2295, R2_n2294, R2_n2293, R2_n2292, R2_n2291, R2_n2290, R2_n2289,
         R2_n2288, R2_n2287, R2_n2286, R2_n2285, R2_n2284, R2_n2283, R2_n2282,
         R2_n2281, R2_n2280, R2_n2279, R2_n2278, R2_n2277, R2_n2276, R2_n2275,
         R2_n2274, R2_n2273, R2_n2272, R2_n2271, R2_n2270, R2_n2269, R2_n2268,
         R2_n2267, R2_n2266, R2_n2265, R2_n2264, R2_n2263, R2_n2262, R2_n2261,
         R2_n2260, R2_n2259, R2_n2258, R2_n2257, R2_n2256, R2_n2255, R2_n2254,
         R2_n2253, R2_n2252, R2_n2251, R2_n2250, R2_n2249, R2_n2248, R2_n2247,
         R2_n2246, R2_n2245, R2_n2244, R2_n2243, R2_n2242, R2_n2241, R2_n2240,
         R2_n2239, R2_n2238, R2_n2237, R2_n2236, R2_n2235, R2_n2234, R2_n2233,
         R2_n2232, R2_n2231, R2_n2230, R2_n2229, R2_n2228, R2_n2227, R2_n2226,
         R2_n2225, R2_n2224, R2_n2223, R2_n2222, R2_n2221, R2_n2220, R2_n2219,
         R2_n2218, R2_n2217, R2_n2216, R2_n2215, R2_n2214, R2_n2213, R2_n2212,
         R2_n2211, R2_n2210, R2_n2209, R2_n2208, R2_n2207, R2_n2206, R2_n2205,
         R2_n2204, R2_n2203, R2_n2202, R2_n2201, R2_n2200, R2_n2199, R2_n2198,
         R2_n2197, R2_n2196, R2_n2195, R2_n2194, R2_n2193, R2_n2192, R2_n2191,
         R2_n2190, R2_n2189, R2_n2188, R2_n2187, R2_n2186, R2_n2185, R2_n2184,
         R2_n2183, R2_n2182, R2_n2181, R2_n2180, R2_n2179, R2_n2178, R2_n2177,
         R2_n2176, R2_n2175, R2_n2174, R2_n2173, R2_n2172, R2_n2171, R2_n2170,
         R2_n2169, R2_n2168, R2_n2167, R2_n2166, R2_n2165, R2_n2164, R2_n2163,
         R2_n2162, R2_n2161, R2_n2160, R2_n2159, R2_n2158, R2_n2157, R2_n2156,
         R2_n2155, R2_n2154, R2_n2153, R2_n2152, R2_n2151, R2_n2150, R2_n2149,
         R2_n2148, R2_n2147, R2_n2146, R2_n2145, R2_n2144, R2_n2143, R2_n2142,
         R2_n2141, R2_n2140, R2_n2139, R2_n2138, R2_n2137, R2_n2136, R2_n2135,
         R2_n2134, R2_n2133, R2_n2132, R2_n2131, R2_n2130, R2_n2129, R2_n2128,
         R2_n2127, R2_n2126, R2_n2125, R2_n2124, R2_n2123, R2_n2122, R2_n2121,
         R2_n2120, R2_n2119, R2_n2118, R2_n2117, R2_n2116, R2_n2115, R2_n2114,
         R2_n2113, R2_n2112, R2_n2111, R2_n2110, R2_n2109, R2_n2108, R2_n2107,
         R2_n2106, R2_n2105, R2_n2104, R2_n2103, R2_n2102, R2_n2101, R2_n2100,
         R2_n2099, R2_n2098, R2_n2097, R2_n2096, R2_n2095, R2_n2094, R2_n2093,
         R2_n2092, R2_n2091, R2_n2090, R2_n2089, R2_n2088, R2_n2087, R2_n2086,
         R2_n2085, R2_n2084, R2_n2083, R2_n2082, R2_n2081, R2_n2080, R2_n2079,
         R2_n2078, R2_n2077, R2_n2076, R2_n2075, R2_n2074, R2_n2073, R2_n2072,
         R2_n2071, R2_n2070, R2_n2069, R2_n2068, R2_n2067, R2_n2066, R2_n2065,
         R2_n2064, R2_n2063, R2_n2062, R2_n2061, R2_n2060, R2_n2059, R2_n2058,
         R2_n2057, R2_n2056, R2_n2055, R2_n2054, R2_n2053, R2_n2052, R2_n2051,
         R2_n2050, R2_n2049, R2_n2048, R2_n2047, R2_n2046, R2_n2045, R2_n2044,
         R2_n2043, R2_n2042, R2_n2041, R2_n2040, R2_n2039, R2_n2038, R2_n2037,
         R2_n2036, R2_n2035, R2_n2034, R2_n2033, R2_n2032, R2_n2031, R2_n2030,
         R2_n2029, R2_n2028, R2_n2027, R2_n2026, R2_n2025, R2_n2024, R2_n2023,
         R2_n2022, R2_n2021, R2_n2020, R2_n2019, R2_n2018, R2_n2017, R2_n2016,
         R2_n2015, R2_n2014, R2_n2013, R2_n2012, R2_n2011, R2_n2010, R2_n2009,
         R2_n2008, R2_n2007, R2_n2006, R2_n2005, R2_n2004, R2_n2003, R2_n2002,
         R2_n2001, R2_n2000, R2_n1999, R2_n1998, R2_n1997, R2_n1996, R2_n1995,
         R2_n1994, R2_n1993, R2_n1992, R2_n1991, R2_n1990, R2_n1989, R2_n1988,
         R2_n1987, R2_n1986, R2_n1985, R2_n1984, R2_n1983, R2_n1982, R2_n1981,
         R2_n1980, R2_n1979, R2_n1978, R2_n1977, R2_n1976, R2_n1975, R2_n1974,
         R2_n1973, R2_n1972, R2_n1971, R2_n1970, R2_n1969, R2_n1968, R2_n1967,
         R2_n1966, R2_n1965, R2_n1964, R2_n1963, R2_n1962, R2_n1961, R2_n1960,
         R2_n1959, R2_n1958, R2_n1957, R2_n1956, R2_n1955, R2_n1954, R2_n1953,
         R2_n1952, R2_n1951, R2_n1950, R2_n1949, R2_n1948, R2_n1947, R2_n1946,
         R2_n1945, R2_n1944, R2_n1943, R2_n1942, R2_n1941, R2_n1940, R2_n1939,
         R2_n1938, R2_n1937, R2_n1936, R2_n1935, R2_n1934, R2_n1933, R2_n1932,
         R2_n1931, R2_n1930, R2_n1929, R2_n1928, R2_n1927, R2_n1926, R2_n1925,
         R2_n1924, R2_n1923, R2_n1922, R2_n1921, R2_n1920, R2_n1919, R2_n1918,
         R2_n1917, R2_n1916, R2_n1915, R2_n1914, R2_n1913, R2_n1912, R2_n1911,
         R2_n1910, R2_n1909, R2_n1908, R2_n1907, R2_n1906, R2_n1905, R2_n1904,
         R2_n1903, R2_n1902, R2_n1901, R2_n1900, R2_n1899, R2_n1898, R2_n1897,
         R2_n1896, R2_n1895, R2_n1894, R2_n1893, R2_n1892, R2_n1891, R2_n1890,
         R2_n1889, R2_n1888, R2_n1887, R2_n1886, R2_n1885, R2_n1884, R2_n1883,
         R2_n1882, R2_n1881, R2_n1880, R2_n1879, R2_n1878, R2_n1877, R2_n1876,
         R2_n1875, R2_n1874, R2_n1873, R2_n1872, R2_n1871, R2_n1870, R2_n1869,
         R2_n1868, R2_n1867, R2_n1866, R2_n1865, R2_n1864, R2_n1863, R2_n1862,
         R2_n1861, R2_n1860, R2_n1859, R2_n1858, R2_n1857, R2_n1856, R2_n1855,
         R2_n1854, R2_n1853, R2_n1852, R2_n1851, R2_n1850, R2_n1849, R2_n1848,
         R2_n1847, R2_n1846, R2_n1845, R2_n1844, R2_n1843, R2_n1842, R2_n1841,
         R2_n1840, R2_n1839, R2_n1838, R2_n1837, R2_n1836, R2_n1835, R2_n1834,
         R2_n1833, R2_n1832, R2_n1831, R2_n1830, R2_n1829, R2_n1828, R2_n1827,
         R2_n1826, R2_n1825, R2_n1824, R2_n1823, R2_n1822, R2_n1821, R2_n1820,
         R2_n1819, R2_n1818, R2_n1817, R2_n1816, R2_n1815, R2_n1814, R2_n1813,
         R2_n1812, R2_n1811, R2_n1810, R2_n1809, R2_n1808, R2_n1807, R2_n1806,
         R2_n1805, R2_n1804, R2_n1802, R2_n1800, R2_n1799, R2_n1798, R2_n1797,
         R2_n1796, R2_n1795, R2_n1794, R2_n1793, R2_n1792, R2_n1791, R2_n1790,
         R2_n1789, R2_n1788, R2_n1787, R2_n1786, R2_n1785, R2_n1784, R2_n1783,
         R2_n1782, R2_n1781, R2_n1780, R2_n1779, R2_n1778, R2_n1777, R2_n1776,
         R2_n1775, R2_n1774, R2_n1773, R2_n1772, R2_n1128, R2_n1127, R2_n1126,
         R2_n1125, R2_n1124, R2_n1123, R2_n1122, R2_n1121, R2_n1120, R2_n1119,
         R2_n1118, R2_n1117, R2_n1116, R2_n1115, R2_n1114, R2_n1113, R2_n1112,
         R2_n1111, R2_n1110, R2_n1109, R2_n1108, R2_n1107, R2_n1106, R2_n1105,
         R2_n1104, R2_n1103, R2_n1102, R2_n1101, R2_n1100, R2_n1099, R2_n1098,
         R2_n1097, R2_n1096, R2_n1095, R2_n1094, R2_n1093, R2_n1092, R2_n1091,
         R2_n1090, R2_n1089, R2_n1088, R2_n1087, R2_n1086, R2_n1085, R2_n1084,
         R2_n1083, R2_n1082, R2_n1081, R2_n1080, R2_n1079, R2_n1078, R2_n1077,
         R2_n1076, R2_n1075, R2_n1074, R2_n1073, R2_n1072, R2_n1071, R2_n1070,
         R2_n1069, R2_n1068, R2_n1067, R2_n1066, R2_n1065, R2_n1064, R2_n1063,
         R2_n1062, R2_n1061, R2_n1060, R2_n1059, R2_n1058, R2_n1057, R2_n1056,
         R2_n1055, R2_n1054, R2_n1053, R2_n1052, R2_n1051, R2_n1050, R2_n1049,
         R2_n1048, R2_n1047, R2_n1046, R2_n1045, R2_n1044, R2_n1043, R2_n1042,
         R2_n1041, R2_n1040, R2_n1039, R2_n1038, R2_n1037, R2_n1036, R2_n1035,
         R2_n1034, R2_n1033, R2_n1032, R2_n1031, R2_n1030, R2_n1029, R2_n1028,
         R2_n1027, R2_n1026, R2_n1025, R2_n1024, R2_n1023, R2_n1022, R2_n1021,
         R2_n1020, R2_n1019, R2_n1018, R2_n1017, R2_n1016, R2_n1015, R2_n1014,
         R2_n1013, R2_n1012, R2_n1011, R2_n1010, R2_n1009, R2_n1008, R2_n1007,
         R2_n1006, R2_n1005, R2_n1004, R2_n1003, R2_n1002, R2_n1001, R2_n614,
         R2_n613, R2_n612, R2_n611, R2_n481, R2_n480, R2_n479, R2_n478,
         R2_n477, R2_n476, R2_n475, R2_n474, R2_n473, R2_n472, R2_n471,
         R2_n470, R2_n469, R2_n468, R2_n467, R2_n466, R2_n465, R2_n464,
         R2_n463, R2_n462, R2_n461, R2_n460, R2_n459, R2_n458, R2_n457,
         R2_n456, R2_n455, R2_n454, R2_n453, R2_n452, R2_n451, R2_n450,
         R2_n449, R2_n448, R2_n447, R2_n446, R2_n445, R2_n444, R2_n443,
         R2_n442, R2_n441, R2_n440, R2_n439, R2_n438, R2_n437, R2_n436,
         R2_n435, R2_n434, R2_n433, R2_n432, R2_n431, R2_n430, R2_n429,
         R2_n428, R2_n427, R2_n426, R2_n425, R2_n424, R2_n423, R2_n422,
         R2_n421, R2_n420, R2_n419, R2_n418, R2_n417, R2_n416, R2_n415,
         R2_n414, R2_n413, R2_n412, R2_n411, R2_n410, R2_n409, R2_n408,
         R2_n407, R2_n406, R2_n405, R2_n404, R2_n403, R2_n402, R2_n401,
         R2_n400, R2_n399, R2_n398, R2_n397, R2_n396, R2_n395, R2_n394,
         R2_n393, R2_n392, R2_n391, R2_n390, R2_n389, R2_n388, R2_n387,
         R2_n386, R2_n385, R2_n384, R2_n383, R2_n382, R2_n381, R2_n380,
         R2_n379, R2_n378, R2_n377, R2_n376, R2_n375, R2_n374, R2_n373,
         R2_n372, R2_n371, R2_n370, R2_n369, R2_n368, R2_n367, R2_n366,
         R2_n365, R2_n364, R2_n363, R2_n362, R2_n361, R2_n360, R2_n359,
         R2_n358, R2_n357, R2_n356, R2_n355, R2_n354, R2_n353, R2_n224,
         R2_n223, R2_n222, R2_n221, R2_n220, R2_n219, R2_n218, R2_n217,
         R2_n216, R2_n215, R2_n214, R2_n213, R2_n212, R2_n211, R2_n210,
         R2_n209, R2_n208, R2_n207, R2_n206, R2_n205, R2_n204, R2_n203,
         R2_n202, R2_n201, R2_n200, R2_n199, R2_n198, R2_n197, R2_n196,
         R2_n195, R2_n194, R2_n193, R2_n192, R2_n191, R2_n190, R2_n189,
         R2_n188, R2_n187, R2_n186, R2_n185, R2_n184, R2_n183, R2_n182,
         R2_n181, R2_n180, R2_n179, R2_n178, R2_n177, R2_n176, R2_n175,
         R2_n174, R2_n173, R2_n172, R2_n171, R2_n170, R2_n169, R2_n168,
         R2_n167, R2_n166, R2_n165, R2_n164, R2_n163, R2_n162, R2_n161,
         R2_n160, R2_n159, R2_n158, R2_n157, R2_n156, R2_n155, R2_n154,
         R2_n153, R2_n152, R2_n151, R2_n150, R2_n149, R2_n148, R2_n147,
         R2_n146, R2_n145, R2_n144, R2_n143, R2_n142, R2_n141, R2_n140,
         R2_n139, R2_n138, R2_n137, R2_n136, R2_n135, R2_n134, R2_n133,
         R2_n132, R2_n131, R2_n129, R2_n128, R2_n127, R2_n126, R2_n125,
         R2_n124, R2_n123, R2_n122, R2_n121, R2_n120, R2_n119, R2_n118,
         R2_n117, R2_n116, R2_n115, R2_n114, R2_n113, R2_n112, R2_n111,
         R2_n110, R2_n109, R2_n108, R2_n107, R2_n106, R2_n105, R2_n104,
         R2_n103, R2_n102, R2_n101, R2_n100, R2_n99, R2_n98, R2_n97, R2_n96,
         R2_n95, R2_n94, R2_n93, R2_n92, R2_n91, R2_n90, R2_n89, R2_n88,
         R2_n87, R2_n86, R2_n85, R2_n84, R2_n83, R2_n82, R2_n81, R2_n80,
         R2_n79, R2_n78, R2_n77, R2_n76, R2_n75, R2_n74, R2_n73, R2_n72,
         R2_n71, R2_n70, R2_n69, R2_n68, R2_n67, R2_n66, R2_n65, R2_n64,
         R2_n63, R2_n62, R2_n61, R2_n60, R2_n59, R2_n58, R2_n57, R2_n56,
         R2_n55, R2_n54, R2_n53, R2_n52, R2_n51, R2_n50, R2_n49, R2_n48,
         R2_n47, R2_n46, R2_n45, R2_n44, R2_n43, R2_n42, R2_n41, R2_n40,
         R2_n39, R2_n38, R2_n37, R2_n36, R2_n35, R2_n34, R2_n33, R2_n32,
         R2_n31, R2_n30, R2_n29, R2_n28, R2_n27, R2_n26, R2_n25, R2_n24,
         R2_n23, R2_n22, R2_n21, R2_n20, R2_n19, R2_n18, R2_n17, R2_n16,
         R2_n15, R2_n14, R2_n13, R2_n12, R2_n11, R2_n10, R2_n9, R2_n8, R2_n7,
         R2_n6, R2_n5, R2_n4, R2_n3, R2_n2, R2_n1, R2_r332_A_3_, R2_r332_A_2_,
         R2_r332_A_1_, R2_r332_A_0_, R2_U16_DATA1_127, R2_U16_DATA1_126,
         R2_U16_DATA1_125, R2_U16_DATA1_124, R2_U16_DATA1_123,
         R2_U16_DATA1_122, R2_U16_DATA1_121, R2_U16_DATA1_120,
         R2_U16_DATA1_119, R2_U16_DATA1_118, R2_U16_DATA1_117,
         R2_U16_DATA1_116, R2_U16_DATA1_115, R2_U16_DATA1_114,
         R2_U16_DATA1_113, R2_U16_DATA1_112, R2_U16_DATA1_111,
         R2_U16_DATA1_110, R2_U16_DATA1_109, R2_U16_DATA1_108,
         R2_U16_DATA1_107, R2_U16_DATA1_106, R2_U16_DATA1_105,
         R2_U16_DATA1_104, R2_U16_DATA1_103, R2_U16_DATA1_102,
         R2_U16_DATA1_101, R2_U16_DATA1_100, R2_U16_DATA1_99, R2_U16_DATA1_98,
         R2_U16_DATA1_97, R2_U16_DATA1_96, R2_U16_DATA1_95, R2_U16_DATA1_94,
         R2_U16_DATA1_93, R2_U16_DATA1_92, R2_U16_DATA1_91, R2_U16_DATA1_90,
         R2_U16_DATA1_89, R2_U16_DATA1_88, R2_U16_DATA1_87, R2_U16_DATA1_86,
         R2_U16_DATA1_85, R2_U16_DATA1_84, R2_U16_DATA1_83, R2_U16_DATA1_82,
         R2_U16_DATA1_81, R2_U16_DATA1_80, R2_U16_DATA1_79, R2_U16_DATA1_78,
         R2_U16_DATA1_77, R2_U16_DATA1_76, R2_U16_DATA1_75, R2_U16_DATA1_74,
         R2_U16_DATA1_73, R2_U16_DATA1_72, R2_U16_DATA1_71, R2_U16_DATA1_70,
         R2_U16_DATA1_69, R2_U16_DATA1_68, R2_U16_DATA1_67, R2_U16_DATA1_66,
         R2_U16_DATA1_65, R2_U16_DATA1_64, R2_U16_DATA1_63, R2_U16_DATA1_62,
         R2_U16_DATA1_61, R2_U16_DATA1_60, R2_U16_DATA1_59, R2_U16_DATA1_58,
         R2_U16_DATA1_57, R2_U16_DATA1_56, R2_U16_DATA1_55, R2_U16_DATA1_54,
         R2_U16_DATA1_53, R2_U16_DATA1_52, R2_U16_DATA1_51, R2_U16_DATA1_50,
         R2_U16_DATA1_49, R2_U16_DATA1_48, R2_U16_DATA1_47, R2_U16_DATA1_46,
         R2_U16_DATA1_45, R2_U16_DATA1_44, R2_U16_DATA1_43, R2_U16_DATA1_42,
         R2_U16_DATA1_41, R2_U16_DATA1_40, R2_U16_DATA1_39, R2_U16_DATA1_38,
         R2_U16_DATA1_37, R2_U16_DATA1_36, R2_U16_DATA1_35, R2_U16_DATA1_34,
         R2_U16_DATA1_33, R2_U16_DATA1_32, R2_U16_DATA1_31, R2_U16_DATA1_30,
         R2_U16_DATA1_29, R2_U16_DATA1_28, R2_U16_DATA1_27, R2_U16_DATA1_26,
         R2_U16_DATA1_25, R2_U16_DATA1_24, R2_U16_DATA1_23, R2_U16_DATA1_22,
         R2_U16_DATA1_21, R2_U16_DATA1_20, R2_U16_DATA1_19, R2_U16_DATA1_18,
         R2_U16_DATA1_17, R2_U16_DATA1_16, R2_U16_DATA1_15, R2_U16_DATA1_14,
         R2_U16_DATA1_13, R2_U16_DATA1_12, R2_U16_DATA1_11, R2_U16_DATA1_10,
         R2_U16_DATA1_9, R2_U16_DATA1_8, R2_U16_DATA1_7, R2_U16_DATA1_6,
         R2_U16_DATA1_5, R2_U16_DATA1_4, R2_U16_DATA1_3, R2_U16_DATA1_2,
         R2_U16_DATA1_1, R2_U16_DATA1_0, R2_U16_DATA2_127, R2_U16_DATA2_126,
         R2_U16_DATA2_125, R2_U16_DATA2_124, R2_U16_DATA2_123,
         R2_U16_DATA2_122, R2_U16_DATA2_121, R2_U16_DATA2_120,
         R2_U16_DATA2_119, R2_U16_DATA2_118, R2_U16_DATA2_117,
         R2_U16_DATA2_116, R2_U16_DATA2_115, R2_U16_DATA2_114,
         R2_U16_DATA2_113, R2_U16_DATA2_112, R2_U16_DATA2_111,
         R2_U16_DATA2_110, R2_U16_DATA2_109, R2_U16_DATA2_108,
         R2_U16_DATA2_107, R2_U16_DATA2_106, R2_U16_DATA2_105,
         R2_U16_DATA2_104, R2_U16_DATA2_103, R2_U16_DATA2_102,
         R2_U16_DATA2_101, R2_U16_DATA2_100, R2_U16_DATA2_99, R2_U16_DATA2_98,
         R2_U16_DATA2_97, R2_U16_DATA2_96, R2_U16_DATA2_95, R2_U16_DATA2_94,
         R2_U16_DATA2_93, R2_U16_DATA2_92, R2_U16_DATA2_91, R2_U16_DATA2_90,
         R2_U16_DATA2_89, R2_U16_DATA2_88, R2_U16_DATA2_87, R2_U16_DATA2_86,
         R2_U16_DATA2_85, R2_U16_DATA2_84, R2_U16_DATA2_83, R2_U16_DATA2_82,
         R2_U16_DATA2_81, R2_U16_DATA2_80, R2_U16_DATA2_79, R2_U16_DATA2_78,
         R2_U16_DATA2_77, R2_U16_DATA2_76, R2_U16_DATA2_75, R2_U16_DATA2_74,
         R2_U16_DATA2_73, R2_U16_DATA2_72, R2_U16_DATA2_71, R2_U16_DATA2_70,
         R2_U16_DATA2_69, R2_U16_DATA2_68, R2_U16_DATA2_67, R2_U16_DATA2_66,
         R2_U16_DATA2_65, R2_U16_DATA2_64, R2_U16_DATA2_63, R2_U16_DATA2_62,
         R2_U16_DATA2_61, R2_U16_DATA2_60, R2_U16_DATA2_59, R2_U16_DATA2_58,
         R2_U16_DATA2_57, R2_U16_DATA2_56, R2_U16_DATA2_55, R2_U16_DATA2_54,
         R2_U16_DATA2_53, R2_U16_DATA2_52, R2_U16_DATA2_51, R2_U16_DATA2_50,
         R2_U16_DATA2_49, R2_U16_DATA2_48, R2_U16_DATA2_47, R2_U16_DATA2_46,
         R2_U16_DATA2_45, R2_U16_DATA2_44, R2_U16_DATA2_43, R2_U16_DATA2_42,
         R2_U16_DATA2_41, R2_U16_DATA2_40, R2_U16_DATA2_39, R2_U16_DATA2_38,
         R2_U16_DATA2_37, R2_U16_DATA2_36, R2_U16_DATA2_35, R2_U16_DATA2_34,
         R2_U16_DATA2_33, R2_U16_DATA2_32, R2_U16_DATA2_31, R2_U16_DATA2_30,
         R2_U16_DATA2_29, R2_U16_DATA2_28, R2_U16_DATA2_27, R2_U16_DATA2_26,
         R2_U16_DATA2_25, R2_U16_DATA2_24, R2_U16_DATA2_23, R2_U16_DATA2_22,
         R2_U16_DATA2_21, R2_U16_DATA2_20, R2_U16_DATA2_19, R2_U16_DATA2_18,
         R2_U16_DATA2_17, R2_U16_DATA2_16, R2_U16_DATA2_15, R2_U16_DATA2_14,
         R2_U16_DATA2_13, R2_U16_DATA2_12, R2_U16_DATA2_11, R2_U16_DATA2_10,
         R2_U16_DATA2_9, R2_U16_DATA2_8, R2_U16_DATA2_7, R2_U16_DATA2_6,
         R2_U16_DATA2_5, R2_U16_DATA2_4, R2_U16_DATA2_3, R2_U16_DATA2_2,
         R2_U16_DATA2_1, R2_U16_DATA2_0, R2_U21_Z_1, R2_U22_Z_1, R2_U23_Z_1,
         R2_U24_Z_1, R2_n1771, R2_n1770, R2_n1769, R2_n1768, R2_n1767,
         R2_n1766, R2_n1765, R2_n1764, R2_n1763, R2_n1762, R2_n1761, R2_n1760,
         R2_n1759, R2_n1758, R2_n1757, R2_n1756, R2_n1755, R2_n1754, R2_n1753,
         R2_n1752, R2_n1751, R2_n1750, R2_n1749, R2_n1748, R2_n1747, R2_n1746,
         R2_n1745, R2_n1744, R2_n1743, R2_n1742, R2_n1741, R2_n1740, R2_n1739,
         R2_n1738, R2_n1737, R2_n1736, R2_n1735, R2_n1734, R2_n1733, R2_n1732,
         R2_n1731, R2_n1730, R2_n1729, R2_n1728, R2_n1727, R2_n1726, R2_n1725,
         R2_n1724, R2_n1723, R2_n1722, R2_n1721, R2_n1720, R2_n1719, R2_n1718,
         R2_n1717, R2_n1716, R2_n1715, R2_n1714, R2_n1713, R2_n1712, R2_n1711,
         R2_n1710, R2_n1709, R2_n1708, R2_n1707, R2_n1706, R2_n1705, R2_n1704,
         R2_n1703, R2_n1702, R2_n1701, R2_n1700, R2_n1699, R2_n1698, R2_n1697,
         R2_n1696, R2_n1695, R2_n1694, R2_n1693, R2_n1692, R2_n1691, R2_n1690,
         R2_n1689, R2_n1688, R2_n1687, R2_n1686, R2_n1685, R2_n1684, R2_n1683,
         R2_n1682, R2_n1681, R2_n1680, R2_n1679, R2_n1678, R2_n1677, R2_n1676,
         R2_n1675, R2_n1674, R2_n1673, R2_n1672, R2_n1671, R2_n1670, R2_n1669,
         R2_n1668, R2_n1667, R2_n1666, R2_n1665, R2_n1664, R2_n1663, R2_n1662,
         R2_n1661, R2_n1660, R2_n1659, R2_n1658, R2_n1657, R2_n1656, R2_n1655,
         R2_n1654, R2_n1653, R2_n1652, R2_n1651, R2_n1650, R2_n1649, R2_n1648,
         R2_n1647, R2_n1646, R2_n1645, R2_n1644, R2_n1643, R2_n1642, R2_n1641,
         R2_n1640, R2_n1639, R2_n1638, R2_n1637, R2_n1636, R2_n1635, R2_n1634,
         R2_n1633, R2_n1632, R2_n1631, R2_n1630, R2_n1629, R2_n1628, R2_n1627,
         R2_n1626, R2_n1625, R2_n1624, R2_n1623, R2_n1622, R2_n1621, R2_n1620,
         R2_n1619, R2_n1618, R2_n1617, R2_n1616, R2_n1615, R2_n1614, R2_n1613,
         R2_n1612, R2_n1611, R2_n1610, R2_n1609, R2_n1608, R2_n1607, R2_n1606,
         R2_n1605, R2_n1604, R2_n1603, R2_n1602, R2_n1601, R2_n1600, R2_n1599,
         R2_n1598, R2_n1597, R2_n1596, R2_n1595, R2_n1594, R2_n1593, R2_n1592,
         R2_n1591, R2_n1590, R2_n1589, R2_n1588, R2_n1587, R2_n1586, R2_n1585,
         R2_n1584, R2_n1583, R2_n1582, R2_n1581, R2_n1580, R2_n1579, R2_n1578,
         R2_n1577, R2_n1576, R2_n1575, R2_n1574, R2_n1573, R2_n1572, R2_n1571,
         R2_n1570, R2_n1569, R2_n1568, R2_n1567, R2_n1566, R2_n1565, R2_n1564,
         R2_n1563, R2_n1562, R2_n1561, R2_n1560, R2_n1559, R2_n1558, R2_n1557,
         R2_n1556, R2_n1555, R2_n1554, R2_n1553, R2_n1552, R2_n1551, R2_n1550,
         R2_n1549, R2_n1548, R2_n1547, R2_n1546, R2_n1545, R2_n1544, R2_n1543,
         R2_n1542, R2_n1541, R2_n1540, R2_n1539, R2_n1538, R2_n1537, R2_n1536,
         R2_n1535, R2_n1534, R2_n1533, R2_n1532, R2_n1531, R2_n1530, R2_n1529,
         R2_n1528, R2_n1527, R2_n1526, R2_n1525, R2_n1524, R2_n1523, R2_n1522,
         R2_n1521, R2_n1520, R2_n1519, R2_n1518, R2_n1517, R2_n1516, R2_n1515,
         R2_n1514, R2_n1513, R2_n1512, R2_n1511, R2_n1510, R2_n1509, R2_n1508,
         R2_n1507, R2_n1506, R2_n1505, R2_n1504, R2_n1503, R2_n1502, R2_n1501,
         R2_n1500, R2_n1499, R2_n1498, R2_n1497, R2_n1496, R2_n1495, R2_n1494,
         R2_n1493, R2_n1492, R2_n1491, R2_n1490, R2_n1489, R2_n1488, R2_n1487,
         R2_n1486, R2_n1485, R2_n1484, R2_n1483, R2_n1482, R2_n1481, R2_n1480,
         R2_n1479, R2_n1478, R2_n1477, R2_n1476, R2_n1475, R2_n1474, R2_n1473,
         R2_n1472, R2_n1471, R2_n1470, R2_n1469, R2_n1468, R2_n1467, R2_n1466,
         R2_n1465, R2_n1464, R2_n1463, R2_n1462, R2_n1461, R2_n1460, R2_n1459,
         R2_n1458, R2_n1457, R2_n1456, R2_n1455, R2_n1454, R2_n1453, R2_n1452,
         R2_n1451, R2_n1450, R2_n1449, R2_n1448, R2_n1447, R2_n1446, R2_n1445,
         R2_n1444, R2_n1443, R2_n1442, R2_n1441, R2_n1440, R2_n1439, R2_n1438,
         R2_n1437, R2_n1436, R2_n1435, R2_n1434, R2_n1433, R2_n1432, R2_n1431,
         R2_n1430, R2_n1429, R2_n1428, R2_n1427, R2_n1426, R2_n1425, R2_n1424,
         R2_n1423, R2_n1422, R2_n1421, R2_n1420, R2_n1419, R2_n1418, R2_n1417,
         R2_n1416, R2_n1415, R2_n1414, R2_n1413, R2_n1412, R2_n1411, R2_n1410,
         R2_n1409, R2_n1408, R2_n1407, R2_n1406, R2_n1405, R2_n1404, R2_n1403,
         R2_n1402, R2_n1401, R2_n1400, R2_n1399, R2_n1398, R2_n1397, R2_n1396,
         R2_n1395, R2_n1394, R2_n1393, R2_n1392, R2_n1391, R2_n1390, R2_n1389,
         R2_n1388, R2_n1387, R2_n1386, R2_n1385, R2_n1384, R2_n1383, R2_n1382,
         R2_n1381, R2_n1380, R2_n1379, R2_n1378, R2_n1377, R2_n1376, R2_n1375,
         R2_n1374, R2_n1373, R2_n1372, R2_n1371, R2_n1370, R2_n1369, R2_n1368,
         R2_n1367, R2_n1366, R2_n1365, R2_n1364, R2_n1363, R2_n1362, R2_n1361,
         R2_n1360, R2_n1359, R2_n1358, R2_n1357, R2_n1356, R2_n1355, R2_n1354,
         R2_n1353, R2_n1352, R2_n1351, R2_n1350, R2_n1349, R2_n1348, R2_n1347,
         R2_n1346, R2_n1345, R2_n1344, R2_n1343, R2_n1342, R2_n1341, R2_n1340,
         R2_n1339, R2_n1338, R2_n1337, R2_n1336, R2_n1335, R2_n1334, R2_n1333,
         R2_n1332, R2_n1331, R2_n1330, R2_n1329, R2_n1328, R2_n1327, R2_n1326,
         R2_n1325, R2_n1324, R2_n1323, R2_n1322, R2_n1321, R2_n1320, R2_n1319,
         R2_n1318, R2_n1317, R2_n1316, R2_n1315, R2_n1314, R2_n1313, R2_n1312,
         R2_n1311, R2_n1310, R2_n1309, R2_n1308, R2_n1307, R2_n1306, R2_n1305,
         R2_n1304, R2_n1303, R2_n1302, R2_n1301, R2_n1300, R2_n1299, R2_n1298,
         R2_n1297, R2_n1296, R2_n1295, R2_n1294, R2_n1293, R2_n1292, R2_n1291,
         R2_n1290, R2_n1289, R2_n1288, R2_n1287, R2_n1286, R2_n1285, R2_n1284,
         R2_n1283, R2_n1282, R2_n1281, R2_n1280, R2_n1279, R2_n1278, R2_n1277,
         R2_n1276, R2_n1275, R2_n1274, R2_n1273, R2_n1272, R2_n1271, R2_n1270,
         R2_n1269, R2_n1268, R2_n1267, R2_n1266, R2_n1265, R2_n1264, R2_n1263,
         R2_n1262, R2_n1261, R2_n1260, R2_n1259, R2_n1258, R2_n1256, R2_n1255,
         R2_n1254, R2_n1253, R2_n1252, R2_n1251, R2_n1250, R2_n1249, R2_n1248,
         R2_n1247, R2_n1246, R2_n1245, R2_n1244, R2_n1243, R2_n1242, R2_n1241,
         R2_n1240, R2_n1239, R2_n1238, R2_n1237, R2_n1236, R2_n1235, R2_n1234,
         R2_n1233, R2_n1232, R2_n1231, R2_n1230, R2_n1229, R2_n1228, R2_n1227,
         R2_n1226, R2_n1225, R2_n1224, R2_n1223, R2_n1222, R2_n1221, R2_n1220,
         R2_n1219, R2_n1218, R2_n1217, R2_n1216, R2_n1215, R2_n1214, R2_n1213,
         R2_n1212, R2_n1211, R2_n1210, R2_n1209, R2_n1208, R2_n1207, R2_n1206,
         R2_n1205, R2_n1204, R2_n1203, R2_n1202, R2_n1201, R2_n1200, R2_n1199,
         R2_n1198, R2_n1197, R2_n1196, R2_n1195, R2_n1194, R2_n1193, R2_n1192,
         R2_n1191, R2_n1190, R2_n1189, R2_n1188, R2_n1187, R2_n1186, R2_n1185,
         R2_n1184, R2_n1183, R2_n1182, R2_n1181, R2_n1180, R2_n1179, R2_n1178,
         R2_n1177, R2_n1176, R2_n1175, R2_n1174, R2_n1173, R2_n1172, R2_n1171,
         R2_n1170, R2_n1169, R2_n1168, R2_n1167, R2_n1166, R2_n1165, R2_n1164,
         R2_n1163, R2_n1162, R2_n1161, R2_n1160, R2_n1159, R2_n1158, R2_n1157,
         R2_n1156, R2_n1155, R2_n1154, R2_n1153, R2_n1152, R2_n1151, R2_n1150,
         R2_n1149, R2_n1148, R2_n1147, R2_n1146, R2_n1145, R2_n1144, R2_n1143,
         R2_n1142, R2_n1141, R2_n1140, R2_n1139, R2_n1138, R2_n1137, R2_n1136,
         R2_n1135, R2_n1134, R2_n1133, R2_n1132, R2_n1131, R2_n1130, R2_n1129,
         R2_n999, R2_n998, R2_n997, R2_n996, R2_n995, R2_n994, R2_n993,
         R2_n992, R2_n991, R2_n990, R2_n989, R2_n988, R2_n987, R2_n986,
         R2_n985, R2_n984, R2_n983, R2_n982, R2_n981, R2_n980, R2_n979,
         R2_n978, R2_n977, R2_n976, R2_n975, R2_n974, R2_n973, R2_n972,
         R2_n971, R2_n970, R2_n969, R2_n968, R2_n967, R2_n966, R2_n965,
         R2_n964, R2_n963, R2_n962, R2_n961, R2_n960, R2_n959, R2_n958,
         R2_n957, R2_n956, R2_n955, R2_n954, R2_n953, R2_n952, R2_n951,
         R2_n950, R2_n949, R2_n948, R2_n947, R2_n946, R2_n945, R2_n944,
         R2_n943, R2_n942, R2_n941, R2_n940, R2_n939, R2_n938, R2_n937,
         R2_n936, R2_n935, R2_n934, R2_n933, R2_n932, R2_n931, R2_n930,
         R2_n929, R2_n928, R2_n927, R2_n926, R2_n925, R2_n924, R2_n923,
         R2_n922, R2_n921, R2_n920, R2_n919, R2_n918, R2_n917, R2_n916,
         R2_n915, R2_n914, R2_n913, R2_n912, R2_n911, R2_n910, R2_n909,
         R2_n908, R2_n907, R2_n906, R2_n905, R2_n904, R2_n903, R2_n902,
         R2_n901, R2_n900, R2_n899, R2_n898, R2_n897, R2_n896, R2_n895,
         R2_n894, R2_n893, R2_n892, R2_n891, R2_n890, R2_n889, R2_n888,
         R2_n887, R2_n886, R2_n885, R2_n884, R2_n883, R2_n882, R2_n881,
         R2_n880, R2_n879, R2_n878, R2_n877, R2_n876, R2_n875, R2_n874,
         R2_n873, R2_n872, R2_n871, R2_n870, R2_n869, R2_n868, R2_n867,
         R2_n866, R2_n865, R2_n864, R2_n863, R2_n862, R2_n861, R2_n860,
         R2_n859, R2_n858, R2_n857, R2_n856, R2_n855, R2_n854, R2_n853,
         R2_n852, R2_n851, R2_n850, R2_n849, R2_n848, R2_n847, R2_n846,
         R2_n845, R2_n844, R2_n843, R2_n842, R2_n841, R2_n840, R2_n839,
         R2_n838, R2_n837, R2_n836, R2_n835, R2_n834, R2_n833, R2_n832,
         R2_n831, R2_n830, R2_n829, R2_n828, R2_n827, R2_n826, R2_n825,
         R2_n824, R2_n823, R2_n822, R2_n821, R2_n820, R2_n819, R2_n818,
         R2_n817, R2_n816, R2_n815, R2_n814, R2_n813, R2_n812, R2_n811,
         R2_n810, R2_n809, R2_n808, R2_n807, R2_n806, R2_n805, R2_n804,
         R2_n803, R2_n802, R2_n801, R2_n800, R2_n799, R2_n798, R2_n797,
         R2_n796, R2_n795, R2_n794, R2_n793, R2_n792, R2_n791, R2_n790,
         R2_n789, R2_n788, R2_n787, R2_n786, R2_n785, R2_n784, R2_n783,
         R2_n782, R2_n781, R2_n780, R2_n779, R2_n778, R2_n777, R2_n776,
         R2_n775, R2_n774, R2_n773, R2_n772, R2_n771, R2_n770, R2_n769,
         R2_n768, R2_n767, R2_n766, R2_n765, R2_n764, R2_n763, R2_n762,
         R2_n761, R2_n760, R2_n759, R2_n758, R2_n757, R2_n756, R2_n755,
         R2_n754, R2_n753, R2_n752, R2_n751, R2_n750, R2_n749, R2_n748,
         R2_n747, R2_n746, R2_n745, R2_n744, R2_n610, R2_n609, R2_n608,
         R2_n607, R2_n606, R2_n605, R2_n604, R2_n603, R2_n602, R2_n601,
         R2_n600, R2_n599, R2_n598, R2_n597, R2_n596, R2_n595, R2_n594,
         R2_n593, R2_n592, R2_n591, R2_n590, R2_n589, R2_n588, R2_n587,
         R2_n586, R2_n585, R2_n584, R2_n583, R2_n582, R2_n581, R2_n580,
         R2_n579, R2_n578, R2_n577, R2_n576, R2_n575, R2_n574, R2_n573,
         R2_n572, R2_n571, R2_n570, R2_n569, R2_n568, R2_n567, R2_n566,
         R2_n565, R2_n564, R2_n563, R2_n562, R2_n561, R2_n560, R2_n559,
         R2_n558, R2_n557, R2_n556, R2_n555, R2_n554, R2_n553, R2_n552,
         R2_n551, R2_n550, R2_n549, R2_n548, R2_n547, R2_n546, R2_n545,
         R2_n544, R2_n543, R2_n542, R2_n541, R2_n540, R2_n539, R2_n538,
         R2_n537, R2_n536, R2_n535, R2_n534, R2_n533, R2_n532, R2_n531,
         R2_n530, R2_n529, R2_n528, R2_n527, R2_n526, R2_n525, R2_n524,
         R2_n523, R2_n522, R2_n521, R2_n520, R2_n519, R2_n518, R2_n517,
         R2_n516, R2_n515, R2_n514, R2_n513, R2_n512, R2_n511, R2_n510,
         R2_n509, R2_n508, R2_n507, R2_n506, R2_n505, R2_n504, R2_n503,
         R2_n502, R2_n501, R2_n500, R2_n499, R2_n498, R2_n497, R2_n496,
         R2_n495, R2_n494, R2_n493, R2_n492, R2_n491, R2_n490, R2_n489,
         R2_n488, R2_n487, R2_n486, R2_n485, R2_n484, R2_n483, R2_n482,
         R2_n352, R2_n351, R2_n350, R2_n349, R2_n348, R2_n347, R2_n346,
         R2_n345, R2_n344, R2_n343, R2_n342, R2_n341, R2_n340, R2_n339,
         R2_n338, R2_n337, R2_n336, R2_n335, R2_n334, R2_n333, R2_n332,
         R2_n331, R2_n330, R2_n329, R2_n328, R2_n327, R2_n326, R2_n325,
         R2_n324, R2_n323, R2_n322, R2_n321, R2_n320, R2_n319, R2_n318,
         R2_n317, R2_n316, R2_n315, R2_n314, R2_n313, R2_n312, R2_n311,
         R2_n310, R2_n309, R2_n308, R2_n307, R2_n306, R2_n305, R2_n304,
         R2_n303, R2_n302, R2_n301, R2_n300, R2_n299, R2_n298, R2_n297,
         R2_n296, R2_n295, R2_n294, R2_n293, R2_n292, R2_n291, R2_n290,
         R2_n289, R2_n288, R2_n287, R2_n286, R2_n285, R2_n284, R2_n283,
         R2_n282, R2_n281, R2_n280, R2_n279, R2_n278, R2_n277, R2_n276,
         R2_n275, R2_n274, R2_n273, R2_n272, R2_n271, R2_n270, R2_n269,
         R2_n268, R2_n267, R2_n266, R2_n265, R2_n264, R2_n263, R2_n262,
         R2_n261, R2_n260, R2_n259, R2_n258, R2_n257, R2_n256, R2_n255,
         R2_n254, R2_n253, R2_n252, R2_n251, R2_n250, R2_n249, R2_n248,
         R2_n247, R2_n246, R2_n245, R2_n244, R2_n243, R2_n242, R2_n241,
         R2_n240, R2_n239, R2_n238, R2_n237, R2_n236, R2_n235, R2_n234,
         R2_n233, R2_n232, R2_n231, R2_n230, R2_n229, R2_n228, R2_n227,
         R2_n226, R2_n225, R2_SB_n629, R2_SB_n628, R2_SB_n627, R2_SB_n626,
         R2_SB_n625, R2_SB_n624, R2_SB_n623, R2_SB_n622, R2_SB_n621,
         R2_SB_n620, R2_SB_n619, R2_SB_n618, R2_SB_n617, R2_SB_n616,
         R2_SB_n615, R2_SB_n614, R2_SB_n572, R2_SB_n571, R2_SB_n570,
         R2_SB_n569, R2_SB_n568, R2_SB_n567, R2_SB_n566, R2_SB_n565,
         R2_SB_n564, R2_SB_n563, R2_SB_n562, R2_SB_n561, R2_SB_n560,
         R2_SB_n559, R2_SB_n558, R2_SB_n557, R2_SB_n556, R2_SB_n555,
         R2_SB_n554, R2_SB_n553, R2_SB_n552, R2_SB_n551, R2_SB_n550,
         R2_SB_n549, R2_SB_n548, R2_SB_n547, R2_SB_n546, R2_SB_n545,
         R2_SB_n544, R2_SB_n543, R2_SB_n542, R2_SB_n541, R2_SB_n540,
         R2_SB_n539, R2_SB_n538, R2_SB_n537, R2_SB_n536, R2_SB_n535,
         R2_SB_n534, R2_SB_n533, R2_SB_n532, R2_SB_n531, R2_SB_n530,
         R2_SB_n529, R2_SB_n528, R2_SB_n527, R2_SB_n526, R2_SB_n525,
         R2_SB_n524, R2_SB_n523, R2_SB_n522, R2_SB_n521, R2_SB_n520,
         R2_SB_n519, R2_SB_n518, R2_SB_n517, R2_SB_n516, R2_SB_n515,
         R2_SB_n514, R2_SB_n513, R2_SB_n512, R2_SB_n511, R2_SB_n510,
         R2_SB_n509, R2_SB_n508, R2_SB_n507, R2_SB_n506, R2_SB_n505,
         R2_SB_n504, R2_SB_n503, R2_SB_n502, R2_SB_n501, R2_SB_n500,
         R2_SB_n499, R2_SB_n498, R2_SB_n497, R2_SB_n496, R2_SB_n495,
         R2_SB_n494, R2_SB_n493, R2_SB_n492, R2_SB_n491, R2_SB_n490,
         R2_SB_n489, R2_SB_n488, R2_SB_n487, R2_SB_n486, R2_SB_n485,
         R2_SB_n484, R2_SB_n483, R2_SB_n482, R2_SB_n481, R2_SB_n480,
         R2_SB_n479, R2_SB_n478, R2_SB_n477, R2_SB_n476, R2_SB_n475,
         R2_SB_n474, R2_SB_n473, R2_SB_n472, R2_SB_n471, R2_SB_n470,
         R2_SB_n469, R2_SB_n468, R2_SB_n467, R2_SB_n466, R2_SB_n465,
         R2_SB_n464, R2_SB_n463, R2_SB_n462, R2_SB_n461, R2_SB_n460,
         R2_SB_n459, R2_SB_n458, R2_SB_n457, R2_SB_n456, R2_SB_n455,
         R2_SB_n454, R2_SB_n453, R2_SB_n452, R2_SB_n451, R2_SB_n450,
         R2_SB_n449, R2_SB_n448, R2_SB_n447, R2_SB_n446, R2_SB_n445,
         R2_SB_n444, R2_SB_n443, R2_SB_n442, R2_SB_n441, R2_SB_n440,
         R2_SB_n439, R2_SB_n438, R2_SB_n437, R2_SB_n436, R2_SB_n435,
         R2_SB_n434, R2_SB_n433, R2_SB_n432, R2_SB_n431, R2_SB_n430,
         R2_SB_n429, R2_SB_n428, R2_SB_n427, R2_SB_n426, R2_SB_n425,
         R2_SB_n424, R2_SB_n423, R2_SB_n422, R2_SB_n421, R2_SB_n420,
         R2_SB_n419, R2_SB_n418, R2_SB_n417, R2_SB_n416, R2_SB_n415,
         R2_SB_n414, R2_SB_n413, R2_SB_n412, R2_SB_n411, R2_SB_n410,
         R2_SB_n409, R2_SB_n408, R2_SB_n407, R2_SB_n406, R2_SB_n405,
         R2_SB_n404, R2_SB_n403, R2_SB_n402, R2_SB_n401, R2_SB_n400,
         R2_SB_n399, R2_SB_n398, R2_SB_n397, R2_SB_n396, R2_SB_n395,
         R2_SB_n394, R2_SB_n393, R2_SB_n392, R2_SB_n391, R2_SB_n390,
         R2_SB_n389, R2_SB_n388, R2_SB_n387, R2_SB_n386, R2_SB_n385,
         R2_SB_n384, R2_SB_n383, R2_SB_n382, R2_SB_n381, R2_SB_n380,
         R2_SB_n379, R2_SB_n378, R2_SB_n377, R2_SB_n376, R2_SB_n375,
         R2_SB_n374, R2_SB_n373, R2_SB_n372, R2_SB_n371, R2_SB_n370,
         R2_SB_n369, R2_SB_n368, R2_SB_n367, R2_SB_n366, R2_SB_n365,
         R2_SB_n364, R2_SB_n363, R2_SB_n362, R2_SB_n361, R2_SB_n360,
         R2_SB_n359, R2_SB_n358, R2_SB_n357, R2_SB_n356, R2_SB_n355,
         R2_SB_n354, R2_SB_n353, R2_SB_n352, R2_SB_n351, R2_SB_n350,
         R2_SB_n349, R2_SB_n348, R2_SB_n347, R2_SB_n346, R2_SB_n345,
         R2_SB_n280, R2_SB_n279, R2_SB_n278, R2_SB_n277, R2_SB_n275,
         R2_SB_n274, R2_SB_n273, R2_SB_n272, R2_SB_n271, R2_SB_n270,
         R2_SB_n269, R2_SB_n268, R2_SB_n267, R2_SB_n266, R2_SB_n265,
         R2_SB_n264, R2_SB_n263, R2_SB_n262, R2_SB_n261, R2_SB_n260,
         R2_SB_n259, R2_SB_n258, R2_SB_n257, R2_SB_n256, R2_SB_n255,
         R2_SB_n254, R2_SB_n253, R2_SB_n252, R2_SB_n251, R2_SB_n250,
         R2_SB_n249, R2_SB_n248, R2_SB_n247, R2_SB_n246, R2_SB_n245,
         R2_SB_n244, R2_SB_n243, R2_SB_n242, R2_SB_n241, R2_SB_n240,
         R2_SB_n239, R2_SB_n238, R2_SB_n237, R2_SB_n236, R2_SB_n235,
         R2_SB_n234, R2_SB_n233, R2_SB_n232, R2_SB_n231, R2_SB_n230,
         R2_SB_n229, R2_SB_n228, R2_SB_n227, R2_SB_n226, R2_SB_n225,
         R2_SB_n224, R2_SB_n223, R2_SB_n222, R2_SB_n221, R2_SB_n220,
         R2_SB_n219, R2_SB_n218, R2_SB_n217, R2_SB_n216, R2_SB_n215,
         R2_SB_n214, R2_SB_n213, R2_SB_n212, R2_SB_n211, R2_SB_n210,
         R2_SB_n209, R2_SB_n208, R2_SB_n207, R2_SB_n206, R2_SB_n205,
         R2_SB_n204, R2_SB_n203, R2_SB_n202, R2_SB_n201, R2_SB_n200,
         R2_SB_n199, R2_SB_n198, R2_SB_n197, R2_SB_n196, R2_SB_n195,
         R2_SB_n194, R2_SB_n193, R2_SB_n192, R2_SB_n191, R2_SB_n190,
         R2_SB_n189, R2_SB_n188, R2_SB_n187, R2_SB_n186, R2_SB_n185,
         R2_SB_n184, R2_SB_n183, R2_SB_n182, R2_SB_n181, R2_SB_n180,
         R2_SB_n179, R2_SB_n178, R2_SB_n177, R2_SB_n48, R2_SB_n47, R2_SB_n46,
         R2_SB_n45, R2_SB_n44, R2_SB_n43, R2_SB_n42, R2_SB_n41, R2_SB_n40,
         R2_SB_n39, R2_SB_n38, R2_SB_n37, R2_SB_n36, R2_SB_n35, R2_SB_n34,
         R2_SB_n33, R2_SB_n32, R2_SB_n31, R2_SB_n30, R2_SB_n29, R2_SB_n28,
         R2_SB_n27, R2_SB_n26, R2_SB_n25, R2_SB_n24, R2_SB_n23, R2_SB_n22,
         R2_SB_n21, R2_SB_n20, R2_SB_n19, R2_SB_n18, R2_SB_n17, R2_SB_n16,
         R2_SB_n15, R2_SB_n14, R2_SB_n13, R2_SB_n12, R2_SB_n11, R2_SB_n10,
         R2_SB_n9, R2_SB_n8, R2_SB_n7, R2_SB_n6, R2_SB_n5, R2_SB_n4, R2_SB_n3,
         R2_SB_n2, R2_SB_n1, R2_SB_add_108_A_3_, R2_SB_add_108_A_2_,
         R2_SB_add_108_A_1_, R2_SB_add_108_A_0_, R2_SB_U4_Z_2, R2_SB_U4_Z_1,
         R2_SB_U4_Z_0, R2_SB_U7_Z_7, R2_SB_U7_Z_6, R2_SB_U7_Z_5, R2_SB_U7_Z_4,
         R2_SB_U7_Z_3, R2_SB_U7_Z_2, R2_SB_U7_Z_1, R2_SB_U7_Z_0, R2_SB_U8_Z_7,
         R2_SB_U8_Z_6, R2_SB_U8_Z_5, R2_SB_U8_Z_4, R2_SB_U8_Z_3, R2_SB_U8_Z_2,
         R2_SB_U8_Z_1, R2_SB_U8_Z_0, R2_SB_U9_Z_7, R2_SB_U9_Z_6, R2_SB_U9_Z_5,
         R2_SB_U9_Z_4, R2_SB_U9_Z_3, R2_SB_U9_Z_2, R2_SB_U9_Z_1, R2_SB_U9_Z_0,
         R2_SB_U10_Z_7, R2_SB_U10_Z_6, R2_SB_U10_Z_5, R2_SB_U10_Z_4,
         R2_SB_U10_Z_3, R2_SB_U10_Z_2, R2_SB_U10_Z_1, R2_SB_U10_Z_0,
         R2_SB_U11_Z_0, R2_SB_n344, R2_SB_n343, R2_SB_n342, R2_SB_n341,
         R2_SB_n340, R2_SB_n339, R2_SB_n338, R2_SB_n337, R2_SB_n336,
         R2_SB_n335, R2_SB_n334, R2_SB_n333, R2_SB_n332, R2_SB_n331,
         R2_SB_n330, R2_SB_n329, R2_SB_n328, R2_SB_n327, R2_SB_n326,
         R2_SB_n325, R2_SB_n324, R2_SB_n323, R2_SB_n322, R2_SB_n321,
         R2_SB_n320, R2_SB_n319, R2_SB_n318, R2_SB_n317, R2_SB_n316,
         R2_SB_n315, R2_SB_n314, R2_SB_n313, R2_SB_n312, R2_SB_n311,
         R2_SB_n310, R2_SB_n309, R2_SB_n308, R2_SB_n307, R2_SB_n306,
         R2_SB_n305, R2_SB_n304, R2_SB_n303, R2_SB_n302, R2_SB_n301,
         R2_SB_n300, R2_SB_n299, R2_SB_n298, R2_SB_n297, R2_SB_n296,
         R2_SB_n295, R2_SB_n294, R2_SB_n293, R2_SB_n292, R2_SB_n291,
         R2_SB_n290, R2_SB_n289, R2_SB_n276, R2_SB_n176, R2_SB_n175,
         R2_SB_n174, R2_SB_n173, R2_SB_n172, R2_SB_n171, R2_SB_n170,
         R2_SB_n169, R2_SB_n168, R2_SB_n167, R2_SB_n166, R2_SB_n165,
         R2_SB_n164, R2_SB_n163, R2_SB_n162, R2_SB_n161, R2_SB_n160,
         R2_SB_n159, R2_SB_n158, R2_SB_n157, R2_SB_n156, R2_SB_n155,
         R2_SB_n154, R2_SB_n153, R2_SB_n152, R2_SB_n151, R2_SB_n150,
         R2_SB_n149, R2_SB_n148, R2_SB_n147, R2_SB_n146, R2_SB_n145,
         R2_SB_n144, R2_SB_n143, R2_SB_n142, R2_SB_n141, R2_SB_n140,
         R2_SB_n139, R2_SB_n138, R2_SB_n137, R2_SB_n136, R2_SB_n135,
         R2_SB_n134, R2_SB_n133, R2_SB_n132, R2_SB_n131, R2_SB_n130,
         R2_SB_n129, R2_SB_n128, R2_SB_n127, R2_SB_n126, R2_SB_n125,
         R2_SB_n124, R2_SB_n123, R2_SB_n122, R2_SB_n121, R2_SB_n120,
         R2_SB_n119, R2_SB_n118, R2_SB_n117, R2_SB_n116, R2_SB_n115,
         R2_SB_n114, R2_SB_n113, R2_SB_n112, R2_SB_n111, R2_SB_n110,
         R2_SB_n109, R2_SB_n108, R2_SB_n107, R2_SB_n106, R2_SB_n105,
         R2_SB_n104, R2_SB_n103, R2_SB_n102, R2_SB_n101, R2_SB_n100, R2_SB_n99,
         R2_SB_n98, R2_SB_n97, R2_SB_n96, R2_SB_n95, R2_SB_n94, R2_SB_n93,
         R2_SB_n92, R2_SB_n91, R2_SB_n90, R2_SB_n89, R2_SB_n88, R2_SB_n87,
         R2_SB_n86, R2_SB_n85, R2_SB_n84, R2_SB_n83, R2_SB_n82, R2_SB_n81,
         R2_SB_n80, R2_SB_n79, R2_SB_n78, R2_SB_n77, R2_SB_n76, R2_SB_n75,
         R2_SB_n74, R2_SB_n73, R2_SB_n72, R2_SB_n71, R2_SB_n70, R2_SB_n69,
         R2_SB_n68, R2_SB_n67, R2_SB_n66, R2_SB_n65, R2_SB_n64, R2_SB_n63,
         R2_SB_n62, R2_SB_n61, R2_SB_n60, R2_SB_n59, R2_SB_n58, R2_SB_n57,
         R2_SB_n56, R2_SB_n55, R2_SB_n54, R2_SB_n53, R2_SB_n52, R2_SB_n51,
         R2_SB_n50, R2_SB_n49, R2_SB_SB1_n911, R2_SB_SB1_n910, R2_SB_SB1_n909,
         R2_SB_SB1_n908, R2_SB_SB1_n907, R2_SB_SB1_n906, R2_SB_SB1_n905,
         R2_SB_SB1_n904, R2_SB_SB1_n903, R2_SB_SB1_n902, R2_SB_SB1_n901,
         R2_SB_SB1_n900, R2_SB_SB1_n899, R2_SB_SB1_n898, R2_SB_SB1_n897,
         R2_SB_SB1_n896, R2_SB_SB1_n895, R2_SB_SB1_n894, R2_SB_SB1_n893,
         R2_SB_SB1_n892, R2_SB_SB1_n891, R2_SB_SB1_n890, R2_SB_SB1_n889,
         R2_SB_SB1_n888, R2_SB_SB1_n887, R2_SB_SB1_n886, R2_SB_SB1_n885,
         R2_SB_SB1_n884, R2_SB_SB1_n883, R2_SB_SB1_n882, R2_SB_SB1_n881,
         R2_SB_SB1_n880, R2_SB_SB1_n879, R2_SB_SB1_n878, R2_SB_SB1_n877,
         R2_SB_SB1_n876, R2_SB_SB1_n875, R2_SB_SB1_n874, R2_SB_SB1_n873,
         R2_SB_SB1_n872, R2_SB_SB1_n871, R2_SB_SB1_n870, R2_SB_SB1_n869,
         R2_SB_SB1_n868, R2_SB_SB1_n867, R2_SB_SB1_n866, R2_SB_SB1_n865,
         R2_SB_SB1_n864, R2_SB_SB1_n863, R2_SB_SB1_n862, R2_SB_SB1_n861,
         R2_SB_SB1_n860, R2_SB_SB1_n859, R2_SB_SB1_n858, R2_SB_SB1_n857,
         R2_SB_SB1_n856, R2_SB_SB1_n855, R2_SB_SB1_n854, R2_SB_SB1_n853,
         R2_SB_SB1_n852, R2_SB_SB1_n851, R2_SB_SB1_n850, R2_SB_SB1_n849,
         R2_SB_SB1_n848, R2_SB_SB1_n847, R2_SB_SB1_n846, R2_SB_SB1_n845,
         R2_SB_SB1_n844, R2_SB_SB1_n843, R2_SB_SB1_n842, R2_SB_SB1_n841,
         R2_SB_SB1_n840, R2_SB_SB1_n839, R2_SB_SB1_n838, R2_SB_SB1_n837,
         R2_SB_SB1_n836, R2_SB_SB1_n835, R2_SB_SB1_n834, R2_SB_SB1_n833,
         R2_SB_SB1_n832, R2_SB_SB1_n831, R2_SB_SB1_n830, R2_SB_SB1_n829,
         R2_SB_SB1_n828, R2_SB_SB1_n827, R2_SB_SB1_n826, R2_SB_SB1_n825,
         R2_SB_SB1_n824, R2_SB_SB1_n823, R2_SB_SB1_n822, R2_SB_SB1_n821,
         R2_SB_SB1_n820, R2_SB_SB1_n819, R2_SB_SB1_n818, R2_SB_SB1_n817,
         R2_SB_SB1_n816, R2_SB_SB1_n815, R2_SB_SB1_n814, R2_SB_SB1_n813,
         R2_SB_SB1_n812, R2_SB_SB1_n811, R2_SB_SB1_n810, R2_SB_SB1_n809,
         R2_SB_SB1_n808, R2_SB_SB1_n807, R2_SB_SB1_n806, R2_SB_SB1_n805,
         R2_SB_SB1_n804, R2_SB_SB1_n803, R2_SB_SB1_n802, R2_SB_SB1_n801,
         R2_SB_SB1_n800, R2_SB_SB1_n799, R2_SB_SB1_n798, R2_SB_SB1_n797,
         R2_SB_SB1_n796, R2_SB_SB1_n795, R2_SB_SB1_n794, R2_SB_SB1_n793,
         R2_SB_SB1_n792, R2_SB_SB1_n791, R2_SB_SB1_n790, R2_SB_SB1_n789,
         R2_SB_SB1_n788, R2_SB_SB1_n787, R2_SB_SB1_n786, R2_SB_SB1_n785,
         R2_SB_SB1_n784, R2_SB_SB1_n783, R2_SB_SB1_n782, R2_SB_SB1_n781,
         R2_SB_SB1_n780, R2_SB_SB1_n779, R2_SB_SB1_n778, R2_SB_SB1_n777,
         R2_SB_SB1_n776, R2_SB_SB1_n775, R2_SB_SB1_n774, R2_SB_SB1_n773,
         R2_SB_SB1_n772, R2_SB_SB1_n771, R2_SB_SB1_n770, R2_SB_SB1_n769,
         R2_SB_SB1_n768, R2_SB_SB1_n767, R2_SB_SB1_n766, R2_SB_SB1_n765,
         R2_SB_SB1_n764, R2_SB_SB1_n763, R2_SB_SB1_n762, R2_SB_SB1_n761,
         R2_SB_SB1_n760, R2_SB_SB1_n759, R2_SB_SB1_n758, R2_SB_SB1_n757,
         R2_SB_SB1_n756, R2_SB_SB1_n755, R2_SB_SB1_n754, R2_SB_SB1_n753,
         R2_SB_SB1_n752, R2_SB_SB1_n751, R2_SB_SB1_n750, R2_SB_SB1_n749,
         R2_SB_SB1_n748, R2_SB_SB1_n747, R2_SB_SB1_n746, R2_SB_SB1_n745,
         R2_SB_SB1_n744, R2_SB_SB1_n743, R2_SB_SB1_n742, R2_SB_SB1_n741,
         R2_SB_SB1_n740, R2_SB_SB1_n739, R2_SB_SB1_n738, R2_SB_SB1_n737,
         R2_SB_SB1_n736, R2_SB_SB1_n735, R2_SB_SB1_n734, R2_SB_SB1_n733,
         R2_SB_SB1_n732, R2_SB_SB1_n731, R2_SB_SB1_n730, R2_SB_SB1_n729,
         R2_SB_SB1_n728, R2_SB_SB1_n727, R2_SB_SB1_n726, R2_SB_SB1_n725,
         R2_SB_SB1_n724, R2_SB_SB1_n723, R2_SB_SB1_n722, R2_SB_SB1_n721,
         R2_SB_SB1_n720, R2_SB_SB1_n719, R2_SB_SB1_n718, R2_SB_SB1_n717,
         R2_SB_SB1_n716, R2_SB_SB1_n715, R2_SB_SB1_n714, R2_SB_SB1_n713,
         R2_SB_SB1_n712, R2_SB_SB1_n711, R2_SB_SB1_n710, R2_SB_SB1_n709,
         R2_SB_SB1_n708, R2_SB_SB1_n707, R2_SB_SB1_n706, R2_SB_SB1_n705,
         R2_SB_SB1_n704, R2_SB_SB1_n703, R2_SB_SB1_n702, R2_SB_SB1_n701,
         R2_SB_SB1_n700, R2_SB_SB1_n699, R2_SB_SB1_n698, R2_SB_SB1_n697,
         R2_SB_SB1_n696, R2_SB_SB1_n695, R2_SB_SB1_n694, R2_SB_SB1_n693,
         R2_SB_SB1_n692, R2_SB_SB1_n691, R2_SB_SB1_n690, R2_SB_SB1_n689,
         R2_SB_SB1_n688, R2_SB_SB1_n687, R2_SB_SB1_n686, R2_SB_SB1_n685,
         R2_SB_SB1_n684, R2_SB_SB1_n683, R2_SB_SB1_n682, R2_SB_SB1_n681,
         R2_SB_SB1_n680, R2_SB_SB1_n679, R2_SB_SB1_n678, R2_SB_SB1_n677,
         R2_SB_SB1_n676, R2_SB_SB1_n675, R2_SB_SB1_n674, R2_SB_SB1_n673,
         R2_SB_SB1_n672, R2_SB_SB1_n671, R2_SB_SB1_n670, R2_SB_SB1_n669,
         R2_SB_SB1_n668, R2_SB_SB1_n667, R2_SB_SB1_n666, R2_SB_SB1_n665,
         R2_SB_SB1_n664, R2_SB_SB1_n663, R2_SB_SB1_n662, R2_SB_SB1_n661,
         R2_SB_SB1_n660, R2_SB_SB1_n659, R2_SB_SB1_n658, R2_SB_SB1_n657,
         R2_SB_SB1_n656, R2_SB_SB1_n655, R2_SB_SB1_n654, R2_SB_SB1_n653,
         R2_SB_SB1_n652, R2_SB_SB1_n651, R2_SB_SB1_n650, R2_SB_SB1_n649,
         R2_SB_SB1_n648, R2_SB_SB1_n647, R2_SB_SB1_n646, R2_SB_SB1_n645,
         R2_SB_SB1_n644, R2_SB_SB1_n643, R2_SB_SB1_n642, R2_SB_SB1_n641,
         R2_SB_SB1_n640, R2_SB_SB1_n639, R2_SB_SB1_n638, R2_SB_SB1_n637,
         R2_SB_SB1_n636, R2_SB_SB1_n635, R2_SB_SB1_n634, R2_SB_SB1_n633,
         R2_SB_SB1_n632, R2_SB_SB1_n631, R2_SB_SB1_n630, R2_SB_SB1_n629,
         R2_SB_SB1_n628, R2_SB_SB1_n627, R2_SB_SB1_n626, R2_SB_SB1_n625,
         R2_SB_SB1_n624, R2_SB_SB1_n623, R2_SB_SB1_n622, R2_SB_SB1_n621,
         R2_SB_SB1_n620, R2_SB_SB1_n619, R2_SB_SB1_n618, R2_SB_SB1_n617,
         R2_SB_SB1_n616, R2_SB_SB1_n615, R2_SB_SB1_n614, R2_SB_SB1_n613,
         R2_SB_SB1_n612, R2_SB_SB1_n611, R2_SB_SB1_n610, R2_SB_SB1_n609,
         R2_SB_SB1_n608, R2_SB_SB1_n607, R2_SB_SB1_n606, R2_SB_SB1_n605,
         R2_SB_SB1_n604, R2_SB_SB1_n603, R2_SB_SB1_n602, R2_SB_SB1_n601,
         R2_SB_SB1_n600, R2_SB_SB1_n599, R2_SB_SB1_n598, R2_SB_SB1_n597,
         R2_SB_SB1_n596, R2_SB_SB1_n595, R2_SB_SB1_n594, R2_SB_SB1_n593,
         R2_SB_SB1_n592, R2_SB_SB1_n591, R2_SB_SB1_n590, R2_SB_SB1_n589,
         R2_SB_SB1_n588, R2_SB_SB1_n587, R2_SB_SB1_n586, R2_SB_SB1_n585,
         R2_SB_SB1_n584, R2_SB_SB1_n583, R2_SB_SB1_n582, R2_SB_SB1_n581,
         R2_SB_SB1_n580, R2_SB_SB1_n579, R2_SB_SB1_n578, R2_SB_SB1_n577,
         R2_SB_SB1_n576, R2_SB_SB1_n575, R2_SB_SB1_n574, R2_SB_SB1_n573,
         R2_SB_SB1_n572, R2_SB_SB1_n571, R2_SB_SB1_n570, R2_SB_SB1_n569,
         R2_SB_SB1_n568, R2_SB_SB1_n567, R2_SB_SB1_n566, R2_SB_SB1_n565,
         R2_SB_SB1_n564, R2_SB_SB1_n563, R2_SB_SB1_n562, R2_SB_SB1_n561,
         R2_SB_SB1_n560, R2_SB_SB1_n559, R2_SB_SB1_n558, R2_SB_SB1_n557,
         R2_SB_SB1_n556, R2_SB_SB1_n555, R2_SB_SB1_n554, R2_SB_SB1_n553,
         R2_SB_SB1_n552, R2_SB_SB1_n551, R2_SB_SB1_n550, R2_SB_SB1_n549,
         R2_SB_SB1_n548, R2_SB_SB1_n547, R2_SB_SB1_n546, R2_SB_SB1_n545,
         R2_SB_SB1_n544, R2_SB_SB1_n543, R2_SB_SB1_n542, R2_SB_SB1_n541,
         R2_SB_SB1_n540, R2_SB_SB1_n539, R2_SB_SB1_n538, R2_SB_SB1_n537,
         R2_SB_SB1_n536, R2_SB_SB1_n535, R2_SB_SB1_n534, R2_SB_SB1_n533,
         R2_SB_SB1_n532, R2_SB_SB1_n531, R2_SB_SB1_n530, R2_SB_SB1_n529,
         R2_SB_SB1_n528, R2_SB_SB1_n527, R2_SB_SB1_n526, R2_SB_SB1_n525,
         R2_SB_SB1_n524, R2_SB_SB1_n523, R2_SB_SB1_n522, R2_SB_SB1_n521,
         R2_SB_SB1_n520, R2_SB_SB1_n519, R2_SB_SB1_n518, R2_SB_SB1_n517,
         R2_SB_SB1_n516, R2_SB_SB1_n515, R2_SB_SB1_n514, R2_SB_SB1_n513,
         R2_SB_SB1_n512, R2_SB_SB1_n511, R2_SB_SB1_n510, R2_SB_SB1_n509,
         R2_SB_SB1_n508, R2_SB_SB1_n507, R2_SB_SB1_n506, R2_SB_SB1_n505,
         R2_SB_SB1_n504, R2_SB_SB1_n503, R2_SB_SB1_n502, R2_SB_SB1_n501,
         R2_SB_SB1_n500, R2_SB_SB1_n499, R2_SB_SB1_n498, R2_SB_SB1_n497,
         R2_SB_SB1_n496, R2_SB_SB1_n495, R2_SB_SB1_n494, R2_SB_SB1_n493,
         R2_SB_SB1_n492, R2_SB_SB1_n491, R2_SB_SB1_n490, R2_SB_SB1_n489,
         R2_SB_SB1_n488, R2_SB_SB1_n487, R2_SB_SB1_n486, R2_SB_SB1_n485,
         R2_SB_SB1_n484, R2_SB_SB1_n483, R2_SB_SB1_n482, R2_SB_SB1_n481,
         R2_SB_SB1_n480, R2_SB_SB1_n479, R2_SB_SB1_n478, R2_SB_SB1_n477,
         R2_SB_SB1_n476, R2_SB_SB1_n475, R2_SB_SB1_n474, R2_SB_SB1_n473,
         R2_SB_SB1_n472, R2_SB_SB1_n471, R2_SB_SB1_n470, R2_SB_SB1_n469,
         R2_SB_SB1_n468, R2_SB_SB1_n467, R2_SB_SB1_n466, R2_SB_SB1_n465,
         R2_SB_SB1_n464, R2_SB_SB1_n463, R2_SB_SB1_n462, R2_SB_SB1_n461,
         R2_SB_SB1_n460, R2_SB_SB1_n459, R2_SB_SB1_n453, R2_SB_SB1_n452,
         R2_SB_SB1_n89, R2_SB_SB1_n87, R2_SB_SB1_n13, R2_SB_SB2_n911,
         R2_SB_SB2_n910, R2_SB_SB2_n909, R2_SB_SB2_n908, R2_SB_SB2_n907,
         R2_SB_SB2_n906, R2_SB_SB2_n905, R2_SB_SB2_n904, R2_SB_SB2_n903,
         R2_SB_SB2_n902, R2_SB_SB2_n901, R2_SB_SB2_n900, R2_SB_SB2_n899,
         R2_SB_SB2_n898, R2_SB_SB2_n897, R2_SB_SB2_n896, R2_SB_SB2_n895,
         R2_SB_SB2_n894, R2_SB_SB2_n893, R2_SB_SB2_n892, R2_SB_SB2_n891,
         R2_SB_SB2_n890, R2_SB_SB2_n889, R2_SB_SB2_n888, R2_SB_SB2_n887,
         R2_SB_SB2_n886, R2_SB_SB2_n885, R2_SB_SB2_n884, R2_SB_SB2_n883,
         R2_SB_SB2_n882, R2_SB_SB2_n881, R2_SB_SB2_n880, R2_SB_SB2_n879,
         R2_SB_SB2_n878, R2_SB_SB2_n877, R2_SB_SB2_n876, R2_SB_SB2_n875,
         R2_SB_SB2_n874, R2_SB_SB2_n873, R2_SB_SB2_n872, R2_SB_SB2_n871,
         R2_SB_SB2_n870, R2_SB_SB2_n869, R2_SB_SB2_n868, R2_SB_SB2_n867,
         R2_SB_SB2_n866, R2_SB_SB2_n865, R2_SB_SB2_n864, R2_SB_SB2_n863,
         R2_SB_SB2_n862, R2_SB_SB2_n861, R2_SB_SB2_n860, R2_SB_SB2_n859,
         R2_SB_SB2_n858, R2_SB_SB2_n857, R2_SB_SB2_n856, R2_SB_SB2_n855,
         R2_SB_SB2_n854, R2_SB_SB2_n853, R2_SB_SB2_n852, R2_SB_SB2_n851,
         R2_SB_SB2_n850, R2_SB_SB2_n849, R2_SB_SB2_n848, R2_SB_SB2_n847,
         R2_SB_SB2_n846, R2_SB_SB2_n845, R2_SB_SB2_n844, R2_SB_SB2_n843,
         R2_SB_SB2_n842, R2_SB_SB2_n841, R2_SB_SB2_n840, R2_SB_SB2_n839,
         R2_SB_SB2_n838, R2_SB_SB2_n837, R2_SB_SB2_n836, R2_SB_SB2_n835,
         R2_SB_SB2_n834, R2_SB_SB2_n833, R2_SB_SB2_n832, R2_SB_SB2_n831,
         R2_SB_SB2_n830, R2_SB_SB2_n829, R2_SB_SB2_n828, R2_SB_SB2_n827,
         R2_SB_SB2_n826, R2_SB_SB2_n825, R2_SB_SB2_n824, R2_SB_SB2_n823,
         R2_SB_SB2_n822, R2_SB_SB2_n821, R2_SB_SB2_n820, R2_SB_SB2_n819,
         R2_SB_SB2_n818, R2_SB_SB2_n817, R2_SB_SB2_n816, R2_SB_SB2_n815,
         R2_SB_SB2_n814, R2_SB_SB2_n813, R2_SB_SB2_n812, R2_SB_SB2_n811,
         R2_SB_SB2_n810, R2_SB_SB2_n809, R2_SB_SB2_n808, R2_SB_SB2_n807,
         R2_SB_SB2_n806, R2_SB_SB2_n805, R2_SB_SB2_n804, R2_SB_SB2_n803,
         R2_SB_SB2_n802, R2_SB_SB2_n801, R2_SB_SB2_n800, R2_SB_SB2_n799,
         R2_SB_SB2_n798, R2_SB_SB2_n797, R2_SB_SB2_n796, R2_SB_SB2_n795,
         R2_SB_SB2_n794, R2_SB_SB2_n793, R2_SB_SB2_n792, R2_SB_SB2_n791,
         R2_SB_SB2_n790, R2_SB_SB2_n789, R2_SB_SB2_n788, R2_SB_SB2_n787,
         R2_SB_SB2_n786, R2_SB_SB2_n785, R2_SB_SB2_n784, R2_SB_SB2_n783,
         R2_SB_SB2_n782, R2_SB_SB2_n781, R2_SB_SB2_n780, R2_SB_SB2_n779,
         R2_SB_SB2_n778, R2_SB_SB2_n777, R2_SB_SB2_n776, R2_SB_SB2_n775,
         R2_SB_SB2_n774, R2_SB_SB2_n773, R2_SB_SB2_n772, R2_SB_SB2_n771,
         R2_SB_SB2_n770, R2_SB_SB2_n769, R2_SB_SB2_n768, R2_SB_SB2_n767,
         R2_SB_SB2_n766, R2_SB_SB2_n765, R2_SB_SB2_n764, R2_SB_SB2_n763,
         R2_SB_SB2_n762, R2_SB_SB2_n761, R2_SB_SB2_n760, R2_SB_SB2_n759,
         R2_SB_SB2_n758, R2_SB_SB2_n757, R2_SB_SB2_n756, R2_SB_SB2_n755,
         R2_SB_SB2_n754, R2_SB_SB2_n753, R2_SB_SB2_n752, R2_SB_SB2_n751,
         R2_SB_SB2_n750, R2_SB_SB2_n749, R2_SB_SB2_n748, R2_SB_SB2_n747,
         R2_SB_SB2_n746, R2_SB_SB2_n745, R2_SB_SB2_n744, R2_SB_SB2_n743,
         R2_SB_SB2_n742, R2_SB_SB2_n741, R2_SB_SB2_n740, R2_SB_SB2_n739,
         R2_SB_SB2_n738, R2_SB_SB2_n737, R2_SB_SB2_n736, R2_SB_SB2_n735,
         R2_SB_SB2_n734, R2_SB_SB2_n733, R2_SB_SB2_n732, R2_SB_SB2_n731,
         R2_SB_SB2_n730, R2_SB_SB2_n729, R2_SB_SB2_n728, R2_SB_SB2_n727,
         R2_SB_SB2_n726, R2_SB_SB2_n725, R2_SB_SB2_n724, R2_SB_SB2_n723,
         R2_SB_SB2_n722, R2_SB_SB2_n721, R2_SB_SB2_n720, R2_SB_SB2_n719,
         R2_SB_SB2_n718, R2_SB_SB2_n717, R2_SB_SB2_n716, R2_SB_SB2_n715,
         R2_SB_SB2_n714, R2_SB_SB2_n713, R2_SB_SB2_n712, R2_SB_SB2_n711,
         R2_SB_SB2_n710, R2_SB_SB2_n709, R2_SB_SB2_n708, R2_SB_SB2_n707,
         R2_SB_SB2_n706, R2_SB_SB2_n705, R2_SB_SB2_n704, R2_SB_SB2_n703,
         R2_SB_SB2_n702, R2_SB_SB2_n701, R2_SB_SB2_n700, R2_SB_SB2_n699,
         R2_SB_SB2_n698, R2_SB_SB2_n697, R2_SB_SB2_n696, R2_SB_SB2_n695,
         R2_SB_SB2_n694, R2_SB_SB2_n693, R2_SB_SB2_n692, R2_SB_SB2_n691,
         R2_SB_SB2_n690, R2_SB_SB2_n689, R2_SB_SB2_n688, R2_SB_SB2_n687,
         R2_SB_SB2_n686, R2_SB_SB2_n685, R2_SB_SB2_n684, R2_SB_SB2_n683,
         R2_SB_SB2_n682, R2_SB_SB2_n681, R2_SB_SB2_n680, R2_SB_SB2_n679,
         R2_SB_SB2_n678, R2_SB_SB2_n677, R2_SB_SB2_n676, R2_SB_SB2_n675,
         R2_SB_SB2_n674, R2_SB_SB2_n673, R2_SB_SB2_n672, R2_SB_SB2_n671,
         R2_SB_SB2_n670, R2_SB_SB2_n669, R2_SB_SB2_n668, R2_SB_SB2_n667,
         R2_SB_SB2_n666, R2_SB_SB2_n665, R2_SB_SB2_n664, R2_SB_SB2_n663,
         R2_SB_SB2_n662, R2_SB_SB2_n661, R2_SB_SB2_n660, R2_SB_SB2_n659,
         R2_SB_SB2_n658, R2_SB_SB2_n657, R2_SB_SB2_n656, R2_SB_SB2_n655,
         R2_SB_SB2_n654, R2_SB_SB2_n653, R2_SB_SB2_n652, R2_SB_SB2_n651,
         R2_SB_SB2_n650, R2_SB_SB2_n649, R2_SB_SB2_n648, R2_SB_SB2_n647,
         R2_SB_SB2_n646, R2_SB_SB2_n645, R2_SB_SB2_n644, R2_SB_SB2_n643,
         R2_SB_SB2_n642, R2_SB_SB2_n641, R2_SB_SB2_n640, R2_SB_SB2_n639,
         R2_SB_SB2_n638, R2_SB_SB2_n637, R2_SB_SB2_n636, R2_SB_SB2_n635,
         R2_SB_SB2_n634, R2_SB_SB2_n633, R2_SB_SB2_n632, R2_SB_SB2_n631,
         R2_SB_SB2_n630, R2_SB_SB2_n629, R2_SB_SB2_n628, R2_SB_SB2_n627,
         R2_SB_SB2_n626, R2_SB_SB2_n625, R2_SB_SB2_n624, R2_SB_SB2_n623,
         R2_SB_SB2_n622, R2_SB_SB2_n621, R2_SB_SB2_n620, R2_SB_SB2_n619,
         R2_SB_SB2_n618, R2_SB_SB2_n617, R2_SB_SB2_n616, R2_SB_SB2_n615,
         R2_SB_SB2_n614, R2_SB_SB2_n613, R2_SB_SB2_n612, R2_SB_SB2_n611,
         R2_SB_SB2_n610, R2_SB_SB2_n609, R2_SB_SB2_n608, R2_SB_SB2_n607,
         R2_SB_SB2_n606, R2_SB_SB2_n605, R2_SB_SB2_n604, R2_SB_SB2_n603,
         R2_SB_SB2_n602, R2_SB_SB2_n601, R2_SB_SB2_n600, R2_SB_SB2_n599,
         R2_SB_SB2_n598, R2_SB_SB2_n597, R2_SB_SB2_n596, R2_SB_SB2_n595,
         R2_SB_SB2_n594, R2_SB_SB2_n593, R2_SB_SB2_n592, R2_SB_SB2_n591,
         R2_SB_SB2_n590, R2_SB_SB2_n589, R2_SB_SB2_n588, R2_SB_SB2_n587,
         R2_SB_SB2_n586, R2_SB_SB2_n585, R2_SB_SB2_n584, R2_SB_SB2_n583,
         R2_SB_SB2_n582, R2_SB_SB2_n581, R2_SB_SB2_n580, R2_SB_SB2_n579,
         R2_SB_SB2_n578, R2_SB_SB2_n577, R2_SB_SB2_n576, R2_SB_SB2_n575,
         R2_SB_SB2_n574, R2_SB_SB2_n573, R2_SB_SB2_n572, R2_SB_SB2_n571,
         R2_SB_SB2_n570, R2_SB_SB2_n569, R2_SB_SB2_n568, R2_SB_SB2_n567,
         R2_SB_SB2_n566, R2_SB_SB2_n565, R2_SB_SB2_n564, R2_SB_SB2_n563,
         R2_SB_SB2_n562, R2_SB_SB2_n561, R2_SB_SB2_n560, R2_SB_SB2_n559,
         R2_SB_SB2_n558, R2_SB_SB2_n557, R2_SB_SB2_n556, R2_SB_SB2_n555,
         R2_SB_SB2_n554, R2_SB_SB2_n553, R2_SB_SB2_n552, R2_SB_SB2_n551,
         R2_SB_SB2_n550, R2_SB_SB2_n549, R2_SB_SB2_n548, R2_SB_SB2_n547,
         R2_SB_SB2_n546, R2_SB_SB2_n545, R2_SB_SB2_n544, R2_SB_SB2_n543,
         R2_SB_SB2_n542, R2_SB_SB2_n541, R2_SB_SB2_n540, R2_SB_SB2_n539,
         R2_SB_SB2_n538, R2_SB_SB2_n537, R2_SB_SB2_n536, R2_SB_SB2_n535,
         R2_SB_SB2_n534, R2_SB_SB2_n533, R2_SB_SB2_n532, R2_SB_SB2_n531,
         R2_SB_SB2_n530, R2_SB_SB2_n529, R2_SB_SB2_n528, R2_SB_SB2_n527,
         R2_SB_SB2_n526, R2_SB_SB2_n525, R2_SB_SB2_n524, R2_SB_SB2_n523,
         R2_SB_SB2_n522, R2_SB_SB2_n521, R2_SB_SB2_n520, R2_SB_SB2_n519,
         R2_SB_SB2_n518, R2_SB_SB2_n517, R2_SB_SB2_n516, R2_SB_SB2_n515,
         R2_SB_SB2_n514, R2_SB_SB2_n513, R2_SB_SB2_n512, R2_SB_SB2_n511,
         R2_SB_SB2_n510, R2_SB_SB2_n509, R2_SB_SB2_n508, R2_SB_SB2_n507,
         R2_SB_SB2_n506, R2_SB_SB2_n505, R2_SB_SB2_n504, R2_SB_SB2_n503,
         R2_SB_SB2_n502, R2_SB_SB2_n501, R2_SB_SB2_n500, R2_SB_SB2_n499,
         R2_SB_SB2_n498, R2_SB_SB2_n497, R2_SB_SB2_n496, R2_SB_SB2_n495,
         R2_SB_SB2_n494, R2_SB_SB2_n493, R2_SB_SB2_n492, R2_SB_SB2_n491,
         R2_SB_SB2_n490, R2_SB_SB2_n489, R2_SB_SB2_n488, R2_SB_SB2_n487,
         R2_SB_SB2_n486, R2_SB_SB2_n485, R2_SB_SB2_n484, R2_SB_SB2_n483,
         R2_SB_SB2_n482, R2_SB_SB2_n481, R2_SB_SB2_n480, R2_SB_SB2_n479,
         R2_SB_SB2_n478, R2_SB_SB2_n477, R2_SB_SB2_n476, R2_SB_SB2_n475,
         R2_SB_SB2_n474, R2_SB_SB2_n473, R2_SB_SB2_n472, R2_SB_SB2_n471,
         R2_SB_SB2_n470, R2_SB_SB2_n469, R2_SB_SB2_n468, R2_SB_SB2_n467,
         R2_SB_SB2_n466, R2_SB_SB2_n465, R2_SB_SB2_n464, R2_SB_SB2_n463,
         R2_SB_SB2_n462, R2_SB_SB2_n461, R2_SB_SB2_n460, R2_SB_SB2_n459,
         R2_SB_SB2_n453, R2_SB_SB2_n452, R2_SB_SB2_n89, R2_SB_SB2_n87,
         R2_SB_SB2_n13, R2_SB_SB3_n911, R2_SB_SB3_n910, R2_SB_SB3_n909,
         R2_SB_SB3_n908, R2_SB_SB3_n907, R2_SB_SB3_n906, R2_SB_SB3_n905,
         R2_SB_SB3_n904, R2_SB_SB3_n903, R2_SB_SB3_n902, R2_SB_SB3_n901,
         R2_SB_SB3_n900, R2_SB_SB3_n899, R2_SB_SB3_n898, R2_SB_SB3_n897,
         R2_SB_SB3_n896, R2_SB_SB3_n895, R2_SB_SB3_n894, R2_SB_SB3_n893,
         R2_SB_SB3_n892, R2_SB_SB3_n891, R2_SB_SB3_n890, R2_SB_SB3_n889,
         R2_SB_SB3_n888, R2_SB_SB3_n887, R2_SB_SB3_n886, R2_SB_SB3_n885,
         R2_SB_SB3_n884, R2_SB_SB3_n883, R2_SB_SB3_n882, R2_SB_SB3_n881,
         R2_SB_SB3_n880, R2_SB_SB3_n879, R2_SB_SB3_n878, R2_SB_SB3_n877,
         R2_SB_SB3_n876, R2_SB_SB3_n875, R2_SB_SB3_n874, R2_SB_SB3_n873,
         R2_SB_SB3_n872, R2_SB_SB3_n871, R2_SB_SB3_n870, R2_SB_SB3_n869,
         R2_SB_SB3_n868, R2_SB_SB3_n867, R2_SB_SB3_n866, R2_SB_SB3_n865,
         R2_SB_SB3_n864, R2_SB_SB3_n863, R2_SB_SB3_n862, R2_SB_SB3_n861,
         R2_SB_SB3_n860, R2_SB_SB3_n859, R2_SB_SB3_n858, R2_SB_SB3_n857,
         R2_SB_SB3_n856, R2_SB_SB3_n855, R2_SB_SB3_n854, R2_SB_SB3_n853,
         R2_SB_SB3_n852, R2_SB_SB3_n851, R2_SB_SB3_n850, R2_SB_SB3_n849,
         R2_SB_SB3_n848, R2_SB_SB3_n847, R2_SB_SB3_n846, R2_SB_SB3_n845,
         R2_SB_SB3_n844, R2_SB_SB3_n843, R2_SB_SB3_n842, R2_SB_SB3_n841,
         R2_SB_SB3_n840, R2_SB_SB3_n839, R2_SB_SB3_n838, R2_SB_SB3_n837,
         R2_SB_SB3_n836, R2_SB_SB3_n835, R2_SB_SB3_n834, R2_SB_SB3_n833,
         R2_SB_SB3_n832, R2_SB_SB3_n831, R2_SB_SB3_n830, R2_SB_SB3_n829,
         R2_SB_SB3_n828, R2_SB_SB3_n827, R2_SB_SB3_n826, R2_SB_SB3_n825,
         R2_SB_SB3_n824, R2_SB_SB3_n823, R2_SB_SB3_n822, R2_SB_SB3_n821,
         R2_SB_SB3_n820, R2_SB_SB3_n819, R2_SB_SB3_n818, R2_SB_SB3_n817,
         R2_SB_SB3_n816, R2_SB_SB3_n815, R2_SB_SB3_n814, R2_SB_SB3_n813,
         R2_SB_SB3_n812, R2_SB_SB3_n811, R2_SB_SB3_n810, R2_SB_SB3_n809,
         R2_SB_SB3_n808, R2_SB_SB3_n807, R2_SB_SB3_n806, R2_SB_SB3_n805,
         R2_SB_SB3_n804, R2_SB_SB3_n803, R2_SB_SB3_n802, R2_SB_SB3_n801,
         R2_SB_SB3_n800, R2_SB_SB3_n799, R2_SB_SB3_n798, R2_SB_SB3_n797,
         R2_SB_SB3_n796, R2_SB_SB3_n795, R2_SB_SB3_n794, R2_SB_SB3_n793,
         R2_SB_SB3_n792, R2_SB_SB3_n791, R2_SB_SB3_n790, R2_SB_SB3_n789,
         R2_SB_SB3_n788, R2_SB_SB3_n787, R2_SB_SB3_n786, R2_SB_SB3_n785,
         R2_SB_SB3_n784, R2_SB_SB3_n783, R2_SB_SB3_n782, R2_SB_SB3_n781,
         R2_SB_SB3_n780, R2_SB_SB3_n779, R2_SB_SB3_n778, R2_SB_SB3_n777,
         R2_SB_SB3_n776, R2_SB_SB3_n775, R2_SB_SB3_n774, R2_SB_SB3_n773,
         R2_SB_SB3_n772, R2_SB_SB3_n771, R2_SB_SB3_n770, R2_SB_SB3_n769,
         R2_SB_SB3_n768, R2_SB_SB3_n767, R2_SB_SB3_n766, R2_SB_SB3_n765,
         R2_SB_SB3_n764, R2_SB_SB3_n763, R2_SB_SB3_n762, R2_SB_SB3_n761,
         R2_SB_SB3_n760, R2_SB_SB3_n759, R2_SB_SB3_n758, R2_SB_SB3_n757,
         R2_SB_SB3_n756, R2_SB_SB3_n755, R2_SB_SB3_n754, R2_SB_SB3_n753,
         R2_SB_SB3_n752, R2_SB_SB3_n751, R2_SB_SB3_n750, R2_SB_SB3_n749,
         R2_SB_SB3_n748, R2_SB_SB3_n747, R2_SB_SB3_n746, R2_SB_SB3_n745,
         R2_SB_SB3_n744, R2_SB_SB3_n743, R2_SB_SB3_n742, R2_SB_SB3_n741,
         R2_SB_SB3_n740, R2_SB_SB3_n739, R2_SB_SB3_n738, R2_SB_SB3_n737,
         R2_SB_SB3_n736, R2_SB_SB3_n735, R2_SB_SB3_n734, R2_SB_SB3_n733,
         R2_SB_SB3_n732, R2_SB_SB3_n731, R2_SB_SB3_n730, R2_SB_SB3_n729,
         R2_SB_SB3_n728, R2_SB_SB3_n727, R2_SB_SB3_n726, R2_SB_SB3_n725,
         R2_SB_SB3_n724, R2_SB_SB3_n723, R2_SB_SB3_n722, R2_SB_SB3_n721,
         R2_SB_SB3_n720, R2_SB_SB3_n719, R2_SB_SB3_n718, R2_SB_SB3_n717,
         R2_SB_SB3_n716, R2_SB_SB3_n715, R2_SB_SB3_n714, R2_SB_SB3_n713,
         R2_SB_SB3_n712, R2_SB_SB3_n711, R2_SB_SB3_n710, R2_SB_SB3_n709,
         R2_SB_SB3_n708, R2_SB_SB3_n707, R2_SB_SB3_n706, R2_SB_SB3_n705,
         R2_SB_SB3_n704, R2_SB_SB3_n703, R2_SB_SB3_n702, R2_SB_SB3_n701,
         R2_SB_SB3_n700, R2_SB_SB3_n699, R2_SB_SB3_n698, R2_SB_SB3_n697,
         R2_SB_SB3_n696, R2_SB_SB3_n695, R2_SB_SB3_n694, R2_SB_SB3_n693,
         R2_SB_SB3_n692, R2_SB_SB3_n691, R2_SB_SB3_n690, R2_SB_SB3_n689,
         R2_SB_SB3_n688, R2_SB_SB3_n687, R2_SB_SB3_n686, R2_SB_SB3_n685,
         R2_SB_SB3_n684, R2_SB_SB3_n683, R2_SB_SB3_n682, R2_SB_SB3_n681,
         R2_SB_SB3_n680, R2_SB_SB3_n679, R2_SB_SB3_n678, R2_SB_SB3_n677,
         R2_SB_SB3_n676, R2_SB_SB3_n675, R2_SB_SB3_n674, R2_SB_SB3_n673,
         R2_SB_SB3_n672, R2_SB_SB3_n671, R2_SB_SB3_n670, R2_SB_SB3_n669,
         R2_SB_SB3_n668, R2_SB_SB3_n667, R2_SB_SB3_n666, R2_SB_SB3_n665,
         R2_SB_SB3_n664, R2_SB_SB3_n663, R2_SB_SB3_n662, R2_SB_SB3_n661,
         R2_SB_SB3_n660, R2_SB_SB3_n659, R2_SB_SB3_n658, R2_SB_SB3_n657,
         R2_SB_SB3_n656, R2_SB_SB3_n655, R2_SB_SB3_n654, R2_SB_SB3_n653,
         R2_SB_SB3_n652, R2_SB_SB3_n651, R2_SB_SB3_n650, R2_SB_SB3_n649,
         R2_SB_SB3_n648, R2_SB_SB3_n647, R2_SB_SB3_n646, R2_SB_SB3_n645,
         R2_SB_SB3_n644, R2_SB_SB3_n643, R2_SB_SB3_n642, R2_SB_SB3_n641,
         R2_SB_SB3_n640, R2_SB_SB3_n639, R2_SB_SB3_n638, R2_SB_SB3_n637,
         R2_SB_SB3_n636, R2_SB_SB3_n635, R2_SB_SB3_n634, R2_SB_SB3_n633,
         R2_SB_SB3_n632, R2_SB_SB3_n631, R2_SB_SB3_n630, R2_SB_SB3_n629,
         R2_SB_SB3_n628, R2_SB_SB3_n627, R2_SB_SB3_n626, R2_SB_SB3_n625,
         R2_SB_SB3_n624, R2_SB_SB3_n623, R2_SB_SB3_n622, R2_SB_SB3_n621,
         R2_SB_SB3_n620, R2_SB_SB3_n619, R2_SB_SB3_n618, R2_SB_SB3_n617,
         R2_SB_SB3_n616, R2_SB_SB3_n615, R2_SB_SB3_n614, R2_SB_SB3_n613,
         R2_SB_SB3_n612, R2_SB_SB3_n611, R2_SB_SB3_n610, R2_SB_SB3_n609,
         R2_SB_SB3_n608, R2_SB_SB3_n607, R2_SB_SB3_n606, R2_SB_SB3_n605,
         R2_SB_SB3_n604, R2_SB_SB3_n603, R2_SB_SB3_n602, R2_SB_SB3_n601,
         R2_SB_SB3_n600, R2_SB_SB3_n599, R2_SB_SB3_n598, R2_SB_SB3_n597,
         R2_SB_SB3_n596, R2_SB_SB3_n595, R2_SB_SB3_n594, R2_SB_SB3_n593,
         R2_SB_SB3_n592, R2_SB_SB3_n591, R2_SB_SB3_n590, R2_SB_SB3_n589,
         R2_SB_SB3_n588, R2_SB_SB3_n587, R2_SB_SB3_n586, R2_SB_SB3_n585,
         R2_SB_SB3_n584, R2_SB_SB3_n583, R2_SB_SB3_n582, R2_SB_SB3_n581,
         R2_SB_SB3_n580, R2_SB_SB3_n579, R2_SB_SB3_n578, R2_SB_SB3_n577,
         R2_SB_SB3_n576, R2_SB_SB3_n575, R2_SB_SB3_n574, R2_SB_SB3_n573,
         R2_SB_SB3_n572, R2_SB_SB3_n571, R2_SB_SB3_n570, R2_SB_SB3_n569,
         R2_SB_SB3_n568, R2_SB_SB3_n567, R2_SB_SB3_n566, R2_SB_SB3_n565,
         R2_SB_SB3_n564, R2_SB_SB3_n563, R2_SB_SB3_n562, R2_SB_SB3_n561,
         R2_SB_SB3_n560, R2_SB_SB3_n559, R2_SB_SB3_n558, R2_SB_SB3_n557,
         R2_SB_SB3_n556, R2_SB_SB3_n555, R2_SB_SB3_n554, R2_SB_SB3_n553,
         R2_SB_SB3_n552, R2_SB_SB3_n551, R2_SB_SB3_n550, R2_SB_SB3_n549,
         R2_SB_SB3_n548, R2_SB_SB3_n547, R2_SB_SB3_n546, R2_SB_SB3_n545,
         R2_SB_SB3_n544, R2_SB_SB3_n543, R2_SB_SB3_n542, R2_SB_SB3_n541,
         R2_SB_SB3_n540, R2_SB_SB3_n539, R2_SB_SB3_n538, R2_SB_SB3_n537,
         R2_SB_SB3_n536, R2_SB_SB3_n535, R2_SB_SB3_n534, R2_SB_SB3_n533,
         R2_SB_SB3_n532, R2_SB_SB3_n531, R2_SB_SB3_n530, R2_SB_SB3_n529,
         R2_SB_SB3_n528, R2_SB_SB3_n527, R2_SB_SB3_n526, R2_SB_SB3_n525,
         R2_SB_SB3_n524, R2_SB_SB3_n523, R2_SB_SB3_n522, R2_SB_SB3_n521,
         R2_SB_SB3_n520, R2_SB_SB3_n519, R2_SB_SB3_n518, R2_SB_SB3_n517,
         R2_SB_SB3_n516, R2_SB_SB3_n515, R2_SB_SB3_n514, R2_SB_SB3_n513,
         R2_SB_SB3_n512, R2_SB_SB3_n511, R2_SB_SB3_n510, R2_SB_SB3_n509,
         R2_SB_SB3_n508, R2_SB_SB3_n507, R2_SB_SB3_n506, R2_SB_SB3_n505,
         R2_SB_SB3_n504, R2_SB_SB3_n503, R2_SB_SB3_n502, R2_SB_SB3_n501,
         R2_SB_SB3_n500, R2_SB_SB3_n499, R2_SB_SB3_n498, R2_SB_SB3_n497,
         R2_SB_SB3_n496, R2_SB_SB3_n495, R2_SB_SB3_n494, R2_SB_SB3_n493,
         R2_SB_SB3_n492, R2_SB_SB3_n491, R2_SB_SB3_n490, R2_SB_SB3_n489,
         R2_SB_SB3_n488, R2_SB_SB3_n487, R2_SB_SB3_n486, R2_SB_SB3_n485,
         R2_SB_SB3_n484, R2_SB_SB3_n483, R2_SB_SB3_n482, R2_SB_SB3_n481,
         R2_SB_SB3_n480, R2_SB_SB3_n479, R2_SB_SB3_n478, R2_SB_SB3_n477,
         R2_SB_SB3_n476, R2_SB_SB3_n475, R2_SB_SB3_n474, R2_SB_SB3_n473,
         R2_SB_SB3_n472, R2_SB_SB3_n471, R2_SB_SB3_n470, R2_SB_SB3_n469,
         R2_SB_SB3_n468, R2_SB_SB3_n467, R2_SB_SB3_n466, R2_SB_SB3_n465,
         R2_SB_SB3_n464, R2_SB_SB3_n463, R2_SB_SB3_n462, R2_SB_SB3_n461,
         R2_SB_SB3_n460, R2_SB_SB3_n459, R2_SB_SB3_n453, R2_SB_SB3_n452,
         R2_SB_SB3_n89, R2_SB_SB3_n87, R2_SB_SB3_n13, R2_SB_SB4_n911,
         R2_SB_SB4_n910, R2_SB_SB4_n909, R2_SB_SB4_n908, R2_SB_SB4_n907,
         R2_SB_SB4_n906, R2_SB_SB4_n905, R2_SB_SB4_n904, R2_SB_SB4_n903,
         R2_SB_SB4_n902, R2_SB_SB4_n901, R2_SB_SB4_n900, R2_SB_SB4_n899,
         R2_SB_SB4_n898, R2_SB_SB4_n897, R2_SB_SB4_n896, R2_SB_SB4_n895,
         R2_SB_SB4_n894, R2_SB_SB4_n893, R2_SB_SB4_n892, R2_SB_SB4_n891,
         R2_SB_SB4_n890, R2_SB_SB4_n889, R2_SB_SB4_n888, R2_SB_SB4_n887,
         R2_SB_SB4_n886, R2_SB_SB4_n885, R2_SB_SB4_n884, R2_SB_SB4_n883,
         R2_SB_SB4_n882, R2_SB_SB4_n881, R2_SB_SB4_n880, R2_SB_SB4_n879,
         R2_SB_SB4_n878, R2_SB_SB4_n877, R2_SB_SB4_n876, R2_SB_SB4_n875,
         R2_SB_SB4_n874, R2_SB_SB4_n873, R2_SB_SB4_n872, R2_SB_SB4_n871,
         R2_SB_SB4_n870, R2_SB_SB4_n869, R2_SB_SB4_n868, R2_SB_SB4_n867,
         R2_SB_SB4_n866, R2_SB_SB4_n865, R2_SB_SB4_n864, R2_SB_SB4_n863,
         R2_SB_SB4_n862, R2_SB_SB4_n861, R2_SB_SB4_n860, R2_SB_SB4_n859,
         R2_SB_SB4_n858, R2_SB_SB4_n857, R2_SB_SB4_n856, R2_SB_SB4_n855,
         R2_SB_SB4_n854, R2_SB_SB4_n853, R2_SB_SB4_n852, R2_SB_SB4_n851,
         R2_SB_SB4_n850, R2_SB_SB4_n849, R2_SB_SB4_n848, R2_SB_SB4_n847,
         R2_SB_SB4_n846, R2_SB_SB4_n845, R2_SB_SB4_n844, R2_SB_SB4_n843,
         R2_SB_SB4_n842, R2_SB_SB4_n841, R2_SB_SB4_n840, R2_SB_SB4_n839,
         R2_SB_SB4_n838, R2_SB_SB4_n837, R2_SB_SB4_n836, R2_SB_SB4_n835,
         R2_SB_SB4_n834, R2_SB_SB4_n833, R2_SB_SB4_n832, R2_SB_SB4_n831,
         R2_SB_SB4_n830, R2_SB_SB4_n829, R2_SB_SB4_n828, R2_SB_SB4_n827,
         R2_SB_SB4_n826, R2_SB_SB4_n825, R2_SB_SB4_n824, R2_SB_SB4_n823,
         R2_SB_SB4_n822, R2_SB_SB4_n821, R2_SB_SB4_n820, R2_SB_SB4_n819,
         R2_SB_SB4_n818, R2_SB_SB4_n817, R2_SB_SB4_n816, R2_SB_SB4_n815,
         R2_SB_SB4_n814, R2_SB_SB4_n813, R2_SB_SB4_n812, R2_SB_SB4_n811,
         R2_SB_SB4_n810, R2_SB_SB4_n809, R2_SB_SB4_n808, R2_SB_SB4_n807,
         R2_SB_SB4_n806, R2_SB_SB4_n805, R2_SB_SB4_n804, R2_SB_SB4_n803,
         R2_SB_SB4_n802, R2_SB_SB4_n801, R2_SB_SB4_n800, R2_SB_SB4_n799,
         R2_SB_SB4_n798, R2_SB_SB4_n797, R2_SB_SB4_n796, R2_SB_SB4_n795,
         R2_SB_SB4_n794, R2_SB_SB4_n793, R2_SB_SB4_n792, R2_SB_SB4_n791,
         R2_SB_SB4_n790, R2_SB_SB4_n789, R2_SB_SB4_n788, R2_SB_SB4_n787,
         R2_SB_SB4_n786, R2_SB_SB4_n785, R2_SB_SB4_n784, R2_SB_SB4_n783,
         R2_SB_SB4_n782, R2_SB_SB4_n781, R2_SB_SB4_n780, R2_SB_SB4_n779,
         R2_SB_SB4_n778, R2_SB_SB4_n777, R2_SB_SB4_n776, R2_SB_SB4_n775,
         R2_SB_SB4_n774, R2_SB_SB4_n773, R2_SB_SB4_n772, R2_SB_SB4_n771,
         R2_SB_SB4_n770, R2_SB_SB4_n769, R2_SB_SB4_n768, R2_SB_SB4_n767,
         R2_SB_SB4_n766, R2_SB_SB4_n765, R2_SB_SB4_n764, R2_SB_SB4_n763,
         R2_SB_SB4_n762, R2_SB_SB4_n761, R2_SB_SB4_n760, R2_SB_SB4_n759,
         R2_SB_SB4_n758, R2_SB_SB4_n757, R2_SB_SB4_n756, R2_SB_SB4_n755,
         R2_SB_SB4_n754, R2_SB_SB4_n753, R2_SB_SB4_n752, R2_SB_SB4_n751,
         R2_SB_SB4_n750, R2_SB_SB4_n749, R2_SB_SB4_n748, R2_SB_SB4_n747,
         R2_SB_SB4_n746, R2_SB_SB4_n745, R2_SB_SB4_n744, R2_SB_SB4_n743,
         R2_SB_SB4_n742, R2_SB_SB4_n741, R2_SB_SB4_n740, R2_SB_SB4_n739,
         R2_SB_SB4_n738, R2_SB_SB4_n737, R2_SB_SB4_n736, R2_SB_SB4_n735,
         R2_SB_SB4_n734, R2_SB_SB4_n733, R2_SB_SB4_n732, R2_SB_SB4_n731,
         R2_SB_SB4_n730, R2_SB_SB4_n729, R2_SB_SB4_n728, R2_SB_SB4_n727,
         R2_SB_SB4_n726, R2_SB_SB4_n725, R2_SB_SB4_n724, R2_SB_SB4_n723,
         R2_SB_SB4_n722, R2_SB_SB4_n721, R2_SB_SB4_n720, R2_SB_SB4_n719,
         R2_SB_SB4_n718, R2_SB_SB4_n717, R2_SB_SB4_n716, R2_SB_SB4_n715,
         R2_SB_SB4_n714, R2_SB_SB4_n713, R2_SB_SB4_n712, R2_SB_SB4_n711,
         R2_SB_SB4_n710, R2_SB_SB4_n709, R2_SB_SB4_n708, R2_SB_SB4_n707,
         R2_SB_SB4_n706, R2_SB_SB4_n705, R2_SB_SB4_n704, R2_SB_SB4_n703,
         R2_SB_SB4_n702, R2_SB_SB4_n701, R2_SB_SB4_n700, R2_SB_SB4_n699,
         R2_SB_SB4_n698, R2_SB_SB4_n697, R2_SB_SB4_n696, R2_SB_SB4_n695,
         R2_SB_SB4_n694, R2_SB_SB4_n693, R2_SB_SB4_n692, R2_SB_SB4_n691,
         R2_SB_SB4_n690, R2_SB_SB4_n689, R2_SB_SB4_n688, R2_SB_SB4_n687,
         R2_SB_SB4_n686, R2_SB_SB4_n685, R2_SB_SB4_n684, R2_SB_SB4_n683,
         R2_SB_SB4_n682, R2_SB_SB4_n681, R2_SB_SB4_n680, R2_SB_SB4_n679,
         R2_SB_SB4_n678, R2_SB_SB4_n677, R2_SB_SB4_n676, R2_SB_SB4_n675,
         R2_SB_SB4_n674, R2_SB_SB4_n673, R2_SB_SB4_n672, R2_SB_SB4_n671,
         R2_SB_SB4_n670, R2_SB_SB4_n669, R2_SB_SB4_n668, R2_SB_SB4_n667,
         R2_SB_SB4_n666, R2_SB_SB4_n665, R2_SB_SB4_n664, R2_SB_SB4_n663,
         R2_SB_SB4_n662, R2_SB_SB4_n661, R2_SB_SB4_n660, R2_SB_SB4_n659,
         R2_SB_SB4_n658, R2_SB_SB4_n657, R2_SB_SB4_n656, R2_SB_SB4_n655,
         R2_SB_SB4_n654, R2_SB_SB4_n653, R2_SB_SB4_n652, R2_SB_SB4_n651,
         R2_SB_SB4_n650, R2_SB_SB4_n649, R2_SB_SB4_n648, R2_SB_SB4_n647,
         R2_SB_SB4_n646, R2_SB_SB4_n645, R2_SB_SB4_n644, R2_SB_SB4_n643,
         R2_SB_SB4_n642, R2_SB_SB4_n641, R2_SB_SB4_n640, R2_SB_SB4_n639,
         R2_SB_SB4_n638, R2_SB_SB4_n637, R2_SB_SB4_n636, R2_SB_SB4_n635,
         R2_SB_SB4_n634, R2_SB_SB4_n633, R2_SB_SB4_n632, R2_SB_SB4_n631,
         R2_SB_SB4_n630, R2_SB_SB4_n629, R2_SB_SB4_n628, R2_SB_SB4_n627,
         R2_SB_SB4_n626, R2_SB_SB4_n625, R2_SB_SB4_n624, R2_SB_SB4_n623,
         R2_SB_SB4_n622, R2_SB_SB4_n621, R2_SB_SB4_n620, R2_SB_SB4_n619,
         R2_SB_SB4_n618, R2_SB_SB4_n617, R2_SB_SB4_n616, R2_SB_SB4_n615,
         R2_SB_SB4_n614, R2_SB_SB4_n613, R2_SB_SB4_n612, R2_SB_SB4_n611,
         R2_SB_SB4_n610, R2_SB_SB4_n609, R2_SB_SB4_n608, R2_SB_SB4_n607,
         R2_SB_SB4_n606, R2_SB_SB4_n605, R2_SB_SB4_n604, R2_SB_SB4_n603,
         R2_SB_SB4_n602, R2_SB_SB4_n601, R2_SB_SB4_n600, R2_SB_SB4_n599,
         R2_SB_SB4_n598, R2_SB_SB4_n597, R2_SB_SB4_n596, R2_SB_SB4_n595,
         R2_SB_SB4_n594, R2_SB_SB4_n593, R2_SB_SB4_n592, R2_SB_SB4_n591,
         R2_SB_SB4_n590, R2_SB_SB4_n589, R2_SB_SB4_n588, R2_SB_SB4_n587,
         R2_SB_SB4_n586, R2_SB_SB4_n585, R2_SB_SB4_n584, R2_SB_SB4_n583,
         R2_SB_SB4_n582, R2_SB_SB4_n581, R2_SB_SB4_n580, R2_SB_SB4_n579,
         R2_SB_SB4_n578, R2_SB_SB4_n577, R2_SB_SB4_n576, R2_SB_SB4_n575,
         R2_SB_SB4_n574, R2_SB_SB4_n573, R2_SB_SB4_n572, R2_SB_SB4_n571,
         R2_SB_SB4_n570, R2_SB_SB4_n569, R2_SB_SB4_n568, R2_SB_SB4_n567,
         R2_SB_SB4_n566, R2_SB_SB4_n565, R2_SB_SB4_n564, R2_SB_SB4_n563,
         R2_SB_SB4_n562, R2_SB_SB4_n561, R2_SB_SB4_n560, R2_SB_SB4_n559,
         R2_SB_SB4_n558, R2_SB_SB4_n557, R2_SB_SB4_n556, R2_SB_SB4_n555,
         R2_SB_SB4_n554, R2_SB_SB4_n553, R2_SB_SB4_n552, R2_SB_SB4_n551,
         R2_SB_SB4_n550, R2_SB_SB4_n549, R2_SB_SB4_n548, R2_SB_SB4_n547,
         R2_SB_SB4_n546, R2_SB_SB4_n545, R2_SB_SB4_n544, R2_SB_SB4_n543,
         R2_SB_SB4_n542, R2_SB_SB4_n541, R2_SB_SB4_n540, R2_SB_SB4_n539,
         R2_SB_SB4_n538, R2_SB_SB4_n537, R2_SB_SB4_n536, R2_SB_SB4_n535,
         R2_SB_SB4_n534, R2_SB_SB4_n533, R2_SB_SB4_n532, R2_SB_SB4_n531,
         R2_SB_SB4_n530, R2_SB_SB4_n529, R2_SB_SB4_n528, R2_SB_SB4_n527,
         R2_SB_SB4_n526, R2_SB_SB4_n525, R2_SB_SB4_n524, R2_SB_SB4_n523,
         R2_SB_SB4_n522, R2_SB_SB4_n521, R2_SB_SB4_n520, R2_SB_SB4_n519,
         R2_SB_SB4_n518, R2_SB_SB4_n517, R2_SB_SB4_n516, R2_SB_SB4_n515,
         R2_SB_SB4_n514, R2_SB_SB4_n513, R2_SB_SB4_n512, R2_SB_SB4_n511,
         R2_SB_SB4_n510, R2_SB_SB4_n509, R2_SB_SB4_n508, R2_SB_SB4_n507,
         R2_SB_SB4_n506, R2_SB_SB4_n505, R2_SB_SB4_n504, R2_SB_SB4_n503,
         R2_SB_SB4_n502, R2_SB_SB4_n501, R2_SB_SB4_n500, R2_SB_SB4_n499,
         R2_SB_SB4_n498, R2_SB_SB4_n497, R2_SB_SB4_n496, R2_SB_SB4_n495,
         R2_SB_SB4_n494, R2_SB_SB4_n493, R2_SB_SB4_n492, R2_SB_SB4_n491,
         R2_SB_SB4_n490, R2_SB_SB4_n489, R2_SB_SB4_n488, R2_SB_SB4_n487,
         R2_SB_SB4_n486, R2_SB_SB4_n485, R2_SB_SB4_n484, R2_SB_SB4_n483,
         R2_SB_SB4_n482, R2_SB_SB4_n481, R2_SB_SB4_n480, R2_SB_SB4_n479,
         R2_SB_SB4_n478, R2_SB_SB4_n477, R2_SB_SB4_n476, R2_SB_SB4_n475,
         R2_SB_SB4_n474, R2_SB_SB4_n473, R2_SB_SB4_n472, R2_SB_SB4_n471,
         R2_SB_SB4_n470, R2_SB_SB4_n469, R2_SB_SB4_n468, R2_SB_SB4_n467,
         R2_SB_SB4_n466, R2_SB_SB4_n465, R2_SB_SB4_n464, R2_SB_SB4_n463,
         R2_SB_SB4_n462, R2_SB_SB4_n461, R2_SB_SB4_n460, R2_SB_SB4_n459,
         R2_SB_SB4_n453, R2_SB_SB4_n452, R2_SB_SB4_n89, R2_SB_SB4_n87,
         R2_SB_SB4_n13, R2_MC1_n338, R2_MC1_n337, R2_MC1_n336, R2_MC1_n335,
         R2_MC1_n334, R2_MC1_n333, R2_MC1_n332, R2_MC1_n331, R2_MC1_n330,
         R2_MC1_n329, R2_MC1_n328, R2_MC1_n327, R2_MC1_n326, R2_MC1_n325,
         R2_MC1_n324, R2_MC1_n323, R2_MC1_n322, R2_MC1_n321, R2_MC1_n320,
         R2_MC1_n319, R2_MC1_n318, R2_MC1_n317, R2_MC1_n316, R2_MC1_n315,
         R2_MC1_n314, R2_MC1_n313, R2_MC1_n312, R2_MC1_n311, R2_MC1_n310,
         R2_MC1_n309, R2_MC1_n308, R2_MC1_n307, R2_MC1_n306, R2_MC1_n305,
         R2_MC1_n304, R2_MC1_n303, R2_MC1_n302, R2_MC1_n301, R2_MC1_n300,
         R2_MC1_n299, R2_MC1_n298, R2_MC1_n297, R2_MC1_n296, R2_MC1_n295,
         R2_MC1_n294, R2_MC1_n293, R2_MC1_n292, R2_MC1_n291, R2_MC1_n290,
         R2_MC1_n289, R2_MC1_n288, R2_MC1_n287, R2_MC1_n286, R2_MC1_n285,
         R2_MC1_n284, R2_MC1_n283, R2_MC1_n282, R2_MC1_n281, R2_MC1_n280,
         R2_MC1_n279, R2_MC1_n278, R2_MC1_n277, R2_MC1_n276, R2_MC1_n275,
         R2_MC1_n274, R2_MC1_n273, R2_MC1_n272, R2_MC1_n271, R2_MC1_n270,
         R2_MC1_n269, R2_MC1_n268, R2_MC1_n267, R2_MC1_n266, R2_MC1_n265,
         R2_MC1_n264, R2_MC1_n263, R2_MC1_n262, R2_MC1_n261, R2_MC1_n260,
         R2_MC1_n259, R2_MC1_n258, R2_MC1_n257, R2_MC1_n256, R2_MC1_n255,
         R2_MC1_n254, R2_MC1_n253, R2_MC1_n252, R2_MC1_n251, R2_MC1_n250,
         R2_MC1_n249, R2_MC1_n248, R2_MC1_n247, R2_MC1_n246, R2_MC1_n245,
         R2_MC1_n244, R2_MC1_n243, R2_MC1_n242, R2_MC1_n241, R2_MC1_n240,
         R2_MC1_n239, R2_MC1_n238, R2_MC1_n237, R2_MC1_n236, R2_MC1_n235,
         R2_MC1_n234, R2_MC1_n233, R2_MC1_n232, R2_MC1_n231, R2_MC1_n230,
         R2_MC1_n229, R2_MC1_n228, R2_MC1_n227, R2_MC1_n226, R2_MC1_n225,
         R2_MC1_n224, R2_MC1_n223, R2_MC1_n222, R2_MC1_n221, R2_MC1_n220,
         R2_MC1_n219, R2_MC1_n218, R2_MC1_n217, R2_MC1_n216, R2_MC1_n215,
         R2_MC1_n214, R2_MC1_n213, R2_MC1_n212, R2_MC1_n211, R2_MC1_n210,
         R2_MC1_n209, R2_MC1_n208, R2_MC1_n207, R2_MC1_n206, R2_MC1_n205,
         R2_MC1_n204, R2_MC1_n203, R2_MC1_n202, R2_MC1_n201, R2_MC1_n200,
         R2_MC1_n199, R2_MC1_n198, R2_MC1_n197, R2_MC1_n196, R2_MC1_n195,
         R2_MC1_n194, R2_MC1_n193, R2_MC1_n192, R2_MC1_n191, R2_MC1_n190,
         R2_MC1_n189, R2_MC1_n188, R2_MC1_n187, R2_MC1_n186, R2_MC1_n185,
         R2_MC1_n184, R2_MC1_n183, R2_MC1_n182, R2_MC1_n181, R2_MC1_n180,
         R2_MC1_n179, R2_MC1_n178, R2_MC1_n177, R2_MC1_n176, R2_MC1_n175,
         R2_MC1_n174, R2_MC1_n173, R2_MC1_n172, R2_MC1_n171, R2_MC1_n170,
         R2_MC1_n169, R2_MC1_n168, R2_MC1_n167, R2_MC1_n166, R2_MC1_n165,
         R2_MC1_n164, R2_MC1_n163, R2_MC1_n162, R2_MC1_n161, R2_MC1_n160,
         R2_MC1_n159, R2_MC1_n158, R2_MC1_n157, R2_MC1_n156, R2_MC1_n155,
         R2_MC1_n154, R2_MC1_n153, R2_MC1_n152, R2_MC1_n151, R2_MC1_n150,
         R2_MC1_n149, R2_MC1_n148, R2_MC1_n147, R2_MC1_n146, R2_MC1_n145,
         R2_MC1_n144, R2_MC1_n143, R2_MC1_n142, R2_MC1_n141, R2_MC1_n140,
         R2_MC1_n139, R2_MC1_n138, R2_MC1_n137, R2_MC1_n136, R2_MC1_n135,
         R2_MC1_n134, R2_MC1_n133, R2_MC1_n132, R2_MC1_n131, R2_MC1_n130,
         R2_MC1_n129, R2_MC1_n128, R2_MC1_n127, R2_MC1_n126, R2_MC1_n125,
         R2_MC1_n124, R2_MC1_n123, R2_MC1_n122, R2_MC1_n121, R2_MC1_n120,
         R2_MC1_n119, R2_MC1_n118, R2_MC1_n117, R2_MC1_n116, R2_MC1_n115,
         R2_MC1_n114, R2_MC1_n113, R2_MC1_n112, R2_MC1_n111, R2_MC1_n110,
         R2_MC1_n109, R2_MC1_n108, R2_MC1_n107, R2_MC1_n106, R2_MC1_n105,
         R2_MC1_n104, R2_MC1_n103, R2_MC1_n102, R2_MC1_n101, R2_MC1_n100,
         R2_MC1_n99, R2_MC1_n98, R2_MC1_n97, R2_MC1_n96, R2_MC1_n95,
         R2_MC1_n94, R2_MC1_n93, R2_MC1_n92, R2_MC1_n91, R2_MC1_n90,
         R2_MC1_n89, R2_MC1_n88, R2_MC1_n87, R2_MC1_n86, R2_MC1_n85,
         R2_MC1_n84, R2_MC1_n83, R2_MC1_n82, R2_MC1_n81, R2_MC1_n80,
         R2_MC1_n79, R2_MC1_n78, R2_MC1_n77, R2_MC1_n76, R2_MC1_n75,
         R2_MC1_n74, R2_MC1_n73, R2_MC1_n72, R2_MC1_n71, R2_MC1_n70,
         R2_MC1_n69, R2_MC1_n68, R2_MC1_n67, R2_MC1_n66, R2_MC1_n65,
         R2_MC1_n64, R2_MC1_n63, R2_MC1_n62, R2_MC1_n61, R2_MC1_n60,
         R2_MC1_n59, R2_MC1_n58, R2_MC1_n57, R2_MC1_n56, R2_MC1_n55,
         R2_MC1_n54, R2_MC1_n53, R2_MC1_n52, R2_MC1_n51, R2_MC1_n50,
         R2_MC1_n49, R2_MC1_n48, R2_MC1_n47, R2_MC1_n46, R2_MC1_n45,
         R2_MC1_n44, R2_MC1_n43, R2_MC1_n42, R2_MC1_n41, R2_MC1_n40,
         R2_MC1_n39, R2_MC1_n38, R2_MC1_n37, R2_MC1_n36, R2_MC1_n35,
         R2_MC1_n34, R2_MC1_n33, R2_MC1_n32, R2_MC1_n31, R2_MC1_n30,
         R2_MC1_n29, R2_MC1_n28, R2_MC1_n27, R2_MC1_n26, R2_MC1_n25,
         R2_MC1_n24, R2_MC1_n23, R2_MC1_n22, R2_MC1_n21, R2_MC1_n20,
         R2_MC1_n19, R2_MC1_n18, R2_MC1_n17, R2_MC1_n16, R2_MC1_n13,
         R2_MC1_n11, R2_MC1_n7, R2_MC1_n4, R2_MC1_n1, EK0_n569, EK0_n568,
         EK0_n567, EK0_n566, EK0_n565, EK0_n564, EK0_n315, EK0_n314, EK0_n313,
         EK0_n312, EK0_n311, EK0_n310, EK0_n309, EK0_n308, EK0_n307, EK0_n306,
         EK0_n305, EK0_n304, EK0_n303, EK0_n302, EK0_n301, EK0_n300, EK0_n299,
         EK0_n298, EK0_n297, EK0_n296, EK0_n295, EK0_n294, EK0_n293, EK0_n292,
         EK0_n291, EK0_n290, EK0_n289, EK0_n288, EK0_n287, EK0_n277, EK0_n276,
         EK0_n274, EK0_n273, EK0_n272, EK0_n271, EK0_n270, EK0_n269, EK0_n268,
         EK0_n267, EK0_n266, EK0_n265, EK0_n264, EK0_n263, EK0_n262, EK0_n261,
         EK0_n260, EK0_n259, EK0_n258, EK0_n257, EK0_n256, EK0_n255, EK0_n254,
         EK0_n253, EK0_n252, EK0_n251, EK0_n250, EK0_n249, EK0_n248, EK0_n247,
         EK0_n246, EK0_n245, EK0_n244, EK0_n243, EK0_n242, EK0_n241, EK0_n240,
         EK0_n239, EK0_n238, EK0_n237, EK0_n236, EK0_n235, EK0_n234, EK0_n233,
         EK0_n232, EK0_n231, EK0_n230, EK0_n229, EK0_n228, EK0_n227, EK0_n226,
         EK0_n225, EK0_n224, EK0_n222, EK0_n221, EK0_n220, EK0_n219, EK0_n218,
         EK0_n217, EK0_n216, EK0_n215, EK0_n214, EK0_n213, EK0_n212, EK0_n211,
         EK0_n210, EK0_n209, EK0_n208, EK0_n207, EK0_n206, EK0_n205, EK0_n204,
         EK0_n203, EK0_n202, EK0_n201, EK0_n200, EK0_n199, EK0_n198, EK0_n197,
         EK0_n196, EK0_n195, EK0_n186, EK0_n185, EK0_n184, EK0_n183, EK0_n182,
         EK0_n181, EK0_n180, EK0_n179, EK0_n26, EK0_n25, EK0_n24, EK0_n23,
         EK0_n22, EK0_n21, EK0_n20, EK0_n19, EK0_n18, EK0_n17, EK0_n16,
         EK0_n15, EK0_n14, EK0_n13, EK0_n12, EK0_n11, EK0_n10, EK0_n9, EK0_n8,
         EK0_n7, EK0_n6, EK0_n5, EK0_n4, EK0_n3, EK0_n2, EK0_n1,
         EK0_add_99_A_1_, EK0_add_99_A_0_, EK0_U4_Z_1, EK0_U4_Z_0, EK0_U9_Z_7,
         EK0_U9_Z_6, EK0_U9_Z_5, EK0_U9_Z_4, EK0_U9_Z_3, EK0_U9_Z_2,
         EK0_U9_Z_1, EK0_U9_Z_0, EK0_n286, EK0_n285, EK0_n284, EK0_n283,
         EK0_n282, EK0_n281, EK0_n280, EK0_n279, EK0_n278, EK0_n275, EK0_n194,
         EK0_n193, EK0_n192, EK0_n191, EK0_n190, EK0_n189, EK0_n188, EK0_n187,
         EK0_n178, EK0_n177, EK0_n176, EK0_n175, EK0_n174, EK0_n173, EK0_n172,
         EK0_n171, EK0_n170, EK0_n169, EK0_n168, EK0_n167, EK0_n166, EK0_n165,
         EK0_n164, EK0_n163, EK0_n162, EK0_n161, EK0_n160, EK0_n159, EK0_n158,
         EK0_n157, EK0_n156, EK0_n155, EK0_n154, EK0_n153, EK0_n152, EK0_n151,
         EK0_n150, EK0_n149, EK0_n148, EK0_n147, EK0_n146, EK0_n145, EK0_n144,
         EK0_n143, EK0_n142, EK0_n141, EK0_n140, EK0_n139, EK0_n138, EK0_n137,
         EK0_n136, EK0_n135, EK0_n134, EK0_n133, EK0_n132, EK0_n131, EK0_n130,
         EK0_n129, EK0_n128, EK0_n127, EK0_n126, EK0_n125, EK0_n124, EK0_n123,
         EK0_n122, EK0_n121, EK0_n120, EK0_n119, EK0_n118, EK0_n117, EK0_n116,
         EK0_n115, EK0_n114, EK0_n113, EK0_n112, EK0_n111, EK0_n110, EK0_n109,
         EK0_n108, EK0_n107, EK0_n106, EK0_n105, EK0_n104, EK0_n103, EK0_n102,
         EK0_n101, EK0_n100, EK0_n99, EK0_n98, EK0_n97, EK0_n96, EK0_n95,
         EK0_n94, EK0_n93, EK0_n92, EK0_n91, EK0_n90, EK0_n89, EK0_n88,
         EK0_n87, EK0_n86, EK0_n85, EK0_n84, EK0_n83, EK0_n82, EK0_n81,
         EK0_n80, EK0_n79, EK0_n78, EK0_n77, EK0_n76, EK0_n75, EK0_n74,
         EK0_n73, EK0_n72, EK0_n71, EK0_n70, EK0_n69, EK0_n68, EK0_n67,
         EK0_n66, EK0_n65, EK0_n64, EK0_n63, EK0_n62, EK0_n61, EK0_n60,
         EK0_n59, EK0_n58, EK0_n57, EK0_n56, EK0_n55, EK0_n54, EK0_n53,
         EK0_n52, EK0_n51, EK0_n50, EK0_n49, EK0_n48, EK0_n47, EK0_n46,
         EK0_n45, EK0_n44, EK0_n43, EK0_n42, EK0_n41, EK0_n40, EK0_n39,
         EK0_n38, EK0_n37, EK0_n36, EK0_n35, EK0_n34, EK0_n33, EK0_n32,
         EK0_n31, EK0_n30, EK0_n29, EK0_n28, EK0_n27, EK0_SB2_n462,
         EK0_SB2_n461, EK0_SB2_n460, EK0_SB2_n459, EK0_SB2_n453, EK0_SB2_n452,
         EK0_SB2_n89, EK0_SB2_n87, EK0_SB2_n13, EK0_SB2_n458, EK0_SB2_n457,
         EK0_SB2_n456, EK0_SB2_n455, EK0_SB2_n454, EK0_SB2_n451, EK0_SB2_n450,
         EK0_SB2_n449, EK0_SB2_n448, EK0_SB2_n447, EK0_SB2_n446, EK0_SB2_n445,
         EK0_SB2_n444, EK0_SB2_n443, EK0_SB2_n442, EK0_SB2_n441, EK0_SB2_n440,
         EK0_SB2_n439, EK0_SB2_n438, EK0_SB2_n437, EK0_SB2_n436, EK0_SB2_n435,
         EK0_SB2_n434, EK0_SB2_n433, EK0_SB2_n432, EK0_SB2_n431, EK0_SB2_n430,
         EK0_SB2_n429, EK0_SB2_n428, EK0_SB2_n427, EK0_SB2_n426, EK0_SB2_n425,
         EK0_SB2_n424, EK0_SB2_n423, EK0_SB2_n422, EK0_SB2_n421, EK0_SB2_n420,
         EK0_SB2_n419, EK0_SB2_n418, EK0_SB2_n417, EK0_SB2_n416, EK0_SB2_n415,
         EK0_SB2_n414, EK0_SB2_n413, EK0_SB2_n412, EK0_SB2_n411, EK0_SB2_n410,
         EK0_SB2_n409, EK0_SB2_n408, EK0_SB2_n407, EK0_SB2_n406, EK0_SB2_n405,
         EK0_SB2_n404, EK0_SB2_n403, EK0_SB2_n402, EK0_SB2_n401, EK0_SB2_n400,
         EK0_SB2_n399, EK0_SB2_n398, EK0_SB2_n397, EK0_SB2_n396, EK0_SB2_n395,
         EK0_SB2_n394, EK0_SB2_n393, EK0_SB2_n392, EK0_SB2_n391, EK0_SB2_n390,
         EK0_SB2_n389, EK0_SB2_n388, EK0_SB2_n387, EK0_SB2_n386, EK0_SB2_n385,
         EK0_SB2_n384, EK0_SB2_n383, EK0_SB2_n382, EK0_SB2_n381, EK0_SB2_n380,
         EK0_SB2_n379, EK0_SB2_n378, EK0_SB2_n377, EK0_SB2_n376, EK0_SB2_n375,
         EK0_SB2_n374, EK0_SB2_n373, EK0_SB2_n372, EK0_SB2_n371, EK0_SB2_n370,
         EK0_SB2_n369, EK0_SB2_n368, EK0_SB2_n367, EK0_SB2_n366, EK0_SB2_n365,
         EK0_SB2_n364, EK0_SB2_n363, EK0_SB2_n362, EK0_SB2_n361, EK0_SB2_n360,
         EK0_SB2_n359, EK0_SB2_n358, EK0_SB2_n357, EK0_SB2_n356, EK0_SB2_n355,
         EK0_SB2_n354, EK0_SB2_n353, EK0_SB2_n352, EK0_SB2_n351, EK0_SB2_n350,
         EK0_SB2_n349, EK0_SB2_n348, EK0_SB2_n347, EK0_SB2_n346, EK0_SB2_n345,
         EK0_SB2_n344, EK0_SB2_n343, EK0_SB2_n342, EK0_SB2_n341, EK0_SB2_n340,
         EK0_SB2_n339, EK0_SB2_n338, EK0_SB2_n337, EK0_SB2_n336, EK0_SB2_n335,
         EK0_SB2_n334, EK0_SB2_n333, EK0_SB2_n332, EK0_SB2_n331, EK0_SB2_n330,
         EK0_SB2_n329, EK0_SB2_n328, EK0_SB2_n327, EK0_SB2_n326, EK0_SB2_n325,
         EK0_SB2_n324, EK0_SB2_n323, EK0_SB2_n322, EK0_SB2_n321, EK0_SB2_n320,
         EK0_SB2_n319, EK0_SB2_n318, EK0_SB2_n317, EK0_SB2_n316, EK0_SB2_n315,
         EK0_SB2_n314, EK0_SB2_n313, EK0_SB2_n312, EK0_SB2_n311, EK0_SB2_n310,
         EK0_SB2_n309, EK0_SB2_n308, EK0_SB2_n307, EK0_SB2_n306, EK0_SB2_n305,
         EK0_SB2_n304, EK0_SB2_n303, EK0_SB2_n302, EK0_SB2_n301, EK0_SB2_n300,
         EK0_SB2_n299, EK0_SB2_n298, EK0_SB2_n297, EK0_SB2_n296, EK0_SB2_n295,
         EK0_SB2_n294, EK0_SB2_n293, EK0_SB2_n292, EK0_SB2_n291, EK0_SB2_n290,
         EK0_SB2_n289, EK0_SB2_n288, EK0_SB2_n287, EK0_SB2_n286, EK0_SB2_n285,
         EK0_SB2_n284, EK0_SB2_n283, EK0_SB2_n282, EK0_SB2_n281, EK0_SB2_n280,
         EK0_SB2_n279, EK0_SB2_n278, EK0_SB2_n277, EK0_SB2_n276, EK0_SB2_n275,
         EK0_SB2_n274, EK0_SB2_n273, EK0_SB2_n272, EK0_SB2_n271, EK0_SB2_n270,
         EK0_SB2_n269, EK0_SB2_n268, EK0_SB2_n267, EK0_SB2_n266, EK0_SB2_n265,
         EK0_SB2_n264, EK0_SB2_n263, EK0_SB2_n262, EK0_SB2_n261, EK0_SB2_n260,
         EK0_SB2_n259, EK0_SB2_n258, EK0_SB2_n257, EK0_SB2_n256, EK0_SB2_n255,
         EK0_SB2_n254, EK0_SB2_n253, EK0_SB2_n252, EK0_SB2_n251, EK0_SB2_n250,
         EK0_SB2_n249, EK0_SB2_n248, EK0_SB2_n247, EK0_SB2_n246, EK0_SB2_n245,
         EK0_SB2_n244, EK0_SB2_n243, EK0_SB2_n242, EK0_SB2_n241, EK0_SB2_n240,
         EK0_SB2_n239, EK0_SB2_n238, EK0_SB2_n237, EK0_SB2_n236, EK0_SB2_n235,
         EK0_SB2_n234, EK0_SB2_n233, EK0_SB2_n232, EK0_SB2_n231, EK0_SB2_n230,
         EK0_SB2_n229, EK0_SB2_n228, EK0_SB2_n227, EK0_SB2_n226, EK0_SB2_n225,
         EK0_SB2_n224, EK0_SB2_n223, EK0_SB2_n222, EK0_SB2_n221, EK0_SB2_n220,
         EK0_SB2_n219, EK0_SB2_n218, EK0_SB2_n217, EK0_SB2_n216, EK0_SB2_n215,
         EK0_SB2_n214, EK0_SB2_n213, EK0_SB2_n212, EK0_SB2_n211, EK0_SB2_n210,
         EK0_SB2_n209, EK0_SB2_n208, EK0_SB2_n207, EK0_SB2_n206, EK0_SB2_n205,
         EK0_SB2_n204, EK0_SB2_n203, EK0_SB2_n202, EK0_SB2_n201, EK0_SB2_n200,
         EK0_SB2_n199, EK0_SB2_n198, EK0_SB2_n197, EK0_SB2_n196, EK0_SB2_n195,
         EK0_SB2_n194, EK0_SB2_n193, EK0_SB2_n192, EK0_SB2_n191, EK0_SB2_n190,
         EK0_SB2_n189, EK0_SB2_n188, EK0_SB2_n187, EK0_SB2_n186, EK0_SB2_n185,
         EK0_SB2_n184, EK0_SB2_n183, EK0_SB2_n182, EK0_SB2_n181, EK0_SB2_n180,
         EK0_SB2_n179, EK0_SB2_n178, EK0_SB2_n177, EK0_SB2_n176, EK0_SB2_n175,
         EK0_SB2_n174, EK0_SB2_n173, EK0_SB2_n172, EK0_SB2_n171, EK0_SB2_n170,
         EK0_SB2_n169, EK0_SB2_n168, EK0_SB2_n167, EK0_SB2_n166, EK0_SB2_n165,
         EK0_SB2_n164, EK0_SB2_n163, EK0_SB2_n162, EK0_SB2_n161, EK0_SB2_n160,
         EK0_SB2_n159, EK0_SB2_n158, EK0_SB2_n157, EK0_SB2_n156, EK0_SB2_n155,
         EK0_SB2_n154, EK0_SB2_n153, EK0_SB2_n152, EK0_SB2_n151, EK0_SB2_n150,
         EK0_SB2_n149, EK0_SB2_n148, EK0_SB2_n147, EK0_SB2_n146, EK0_SB2_n145,
         EK0_SB2_n144, EK0_SB2_n143, EK0_SB2_n142, EK0_SB2_n141, EK0_SB2_n140,
         EK0_SB2_n139, EK0_SB2_n138, EK0_SB2_n137, EK0_SB2_n136, EK0_SB2_n135,
         EK0_SB2_n134, EK0_SB2_n133, EK0_SB2_n132, EK0_SB2_n131, EK0_SB2_n130,
         EK0_SB2_n129, EK0_SB2_n128, EK0_SB2_n127, EK0_SB2_n126, EK0_SB2_n125,
         EK0_SB2_n124, EK0_SB2_n123, EK0_SB2_n122, EK0_SB2_n121, EK0_SB2_n120,
         EK0_SB2_n119, EK0_SB2_n118, EK0_SB2_n117, EK0_SB2_n116, EK0_SB2_n115,
         EK0_SB2_n114, EK0_SB2_n113, EK0_SB2_n112, EK0_SB2_n111, EK0_SB2_n110,
         EK0_SB2_n109, EK0_SB2_n108, EK0_SB2_n107, EK0_SB2_n106, EK0_SB2_n105,
         EK0_SB2_n104, EK0_SB2_n103, EK0_SB2_n102, EK0_SB2_n101, EK0_SB2_n100,
         EK0_SB2_n99, EK0_SB2_n98, EK0_SB2_n97, EK0_SB2_n96, EK0_SB2_n95,
         EK0_SB2_n94, EK0_SB2_n93, EK0_SB2_n92, EK0_SB2_n91, EK0_SB2_n90,
         EK0_SB2_n88, EK0_SB2_n86, EK0_SB2_n85, EK0_SB2_n84, EK0_SB2_n83,
         EK0_SB2_n82, EK0_SB2_n81, EK0_SB2_n80, EK0_SB2_n79, EK0_SB2_n78,
         EK0_SB2_n77, EK0_SB2_n76, EK0_SB2_n75, EK0_SB2_n74, EK0_SB2_n73,
         EK0_SB2_n72, EK0_SB2_n71, EK0_SB2_n70, EK0_SB2_n69, EK0_SB2_n68,
         EK0_SB2_n67, EK0_SB2_n66, EK0_SB2_n65, EK0_SB2_n64, EK0_SB2_n63,
         EK0_SB2_n62, EK0_SB2_n61, EK0_SB2_n60, EK0_SB2_n59, EK0_SB2_n58,
         EK0_SB2_n57, EK0_SB2_n56, EK0_SB2_n55, EK0_SB2_n54, EK0_SB2_n53,
         EK0_SB2_n52, EK0_SB2_n51, EK0_SB2_n50, EK0_SB2_n49, EK0_SB2_n48,
         EK0_SB2_n47, EK0_SB2_n46, EK0_SB2_n45, EK0_SB2_n44, EK0_SB2_n43,
         EK0_SB2_n42, EK0_SB2_n41, EK0_SB2_n40, EK0_SB2_n39, EK0_SB2_n38,
         EK0_SB2_n37, EK0_SB2_n36, EK0_SB2_n35, EK0_SB2_n34, EK0_SB2_n33,
         EK0_SB2_n32, EK0_SB2_n31, EK0_SB2_n30, EK0_SB2_n29, EK0_SB2_n28,
         EK0_SB2_n27, EK0_SB2_n26, EK0_SB2_n25, EK0_SB2_n24, EK0_SB2_n23,
         EK0_SB2_n22, EK0_SB2_n21, EK0_SB2_n20, EK0_SB2_n19, EK0_SB2_n18,
         EK0_SB2_n17, EK0_SB2_n16, EK0_SB2_n15, EK0_SB2_n14, EK0_SB2_n12,
         EK0_SB2_n11, EK0_SB2_n10, EK0_SB2_n9, EK0_SB2_n8, EK0_SB2_n7,
         EK0_SB2_n6, EK0_SB2_n5, EK0_SB2_n4, EK0_SB2_n3, EK0_SB2_n2,
         EK0_SB2_n1;
  wire   [3124:2997] n;
  wire   [616:743] R2_n;
  wire   [281:288] R2_SB_n;

  DFF_X1 cnt_reg_0_ ( .D(n5407), .CK(clk), .Q(r424_A_0_), .QN(n4599) );
  DLH_X1 round_reg ( .G(n5471), .D(n5408), .Q(n3391) );
  DLH_X1 round_in_data_reg_98_ ( .G(n5471), .D(U49_Z_98), .Q(n3618) );
  DFF_X1 rstR_reg ( .D(n5405), .CK(clk), .Q(n3261) );
  DFF_X1 rstk_reg ( .D(n5405), .CK(clk), .Q(n2995) );
  DFF_X1 ready_reg ( .D(n5402), .CK(clk), .Q(ready), .QN(n4458) );
  DFF_X1 cnt_reg_1_ ( .D(n5403), .CK(clk), .Q(r424_A_1_), .QN(n4598) );
  DFF_X1 cnt_reg_2_ ( .D(n5404), .CK(clk), .Q(r424_A_2_), .QN(n4596) );
  DFF_X1 cnt_reg_3_ ( .D(n5406), .CK(clk), .Q(r424_A_3_), .QN(n4594) );
  DLH_X1 rcon_index_reg_3_ ( .G(n5473), .D(U51_Z_3), .Q(n3128) );
  DLH_X1 rcon_index_reg_2_ ( .G(n5473), .D(U51_Z_2), .Q(n3127) );
  DLH_X1 rcon_index_reg_0_ ( .G(n5474), .D(U51_Z_0), .Q(n3125) );
  DLH_X1 rcon_index_reg_1_ ( .G(n5475), .D(U51_Z_1), .Q(n3126) );
  DFF_X1 expanded_key_reg_127_ ( .D(n4071), .CK(clk), .Q(U99_DATA1_127) );
  DLH_X1 round_in_key_reg_127_ ( .G(n5471), .D(U99_DATA1_127), .Q(n3519) );
  DLH_X1 expanded_key_in_reg_127_ ( .G(n5473), .D(n4330), .Q(n3260) );
  DFF_X1 expanded_key_reg_0_ ( .D(n4170), .CK(clk), .Q(U99_DATA1_0) );
  DLH_X1 round_in_key_reg_0_ ( .G(n5471), .D(U99_DATA1_0), .Q(n3392) );
  DLH_X1 expanded_key_in_reg_0_ ( .G(n5472), .D(n4457), .Q(n3133) );
  DFF_X1 expanded_key_reg_1_ ( .D(n4169), .CK(clk), .Q(U99_DATA1_1) );
  DLH_X1 round_in_key_reg_1_ ( .G(n5470), .D(U99_DATA1_1), .Q(n3393) );
  DLH_X1 expanded_key_in_reg_1_ ( .G(n5472), .D(n4456), .Q(n3134) );
  DFF_X1 expanded_key_reg_2_ ( .D(n4168), .CK(clk), .Q(U99_DATA1_2) );
  DLH_X1 round_in_key_reg_2_ ( .G(n5470), .D(U99_DATA1_2), .Q(n3394) );
  DLH_X1 expanded_key_in_reg_2_ ( .G(U47_Z_1), .D(n4455), .Q(n3135) );
  DFF_X1 expanded_key_reg_3_ ( .D(n4167), .CK(clk), .Q(U99_DATA1_3) );
  DLH_X1 round_in_key_reg_3_ ( .G(n5470), .D(U99_DATA1_3), .Q(n3395) );
  DLH_X1 expanded_key_in_reg_3_ ( .G(n5472), .D(n4454), .Q(n3136) );
  DFF_X1 expanded_key_reg_4_ ( .D(n4166), .CK(clk), .Q(U99_DATA1_4) );
  DLH_X1 round_in_key_reg_4_ ( .G(n5470), .D(U99_DATA1_4), .Q(n3396) );
  DLH_X1 expanded_key_in_reg_4_ ( .G(n5473), .D(n4453), .Q(n3137) );
  DFF_X1 expanded_key_reg_5_ ( .D(n4165), .CK(clk), .Q(U99_DATA1_5) );
  DLH_X1 round_in_key_reg_5_ ( .G(n5470), .D(U99_DATA1_5), .Q(n3397) );
  DLH_X1 expanded_key_in_reg_5_ ( .G(n5474), .D(n4452), .Q(n3138) );
  DFF_X1 expanded_key_reg_6_ ( .D(n4164), .CK(clk), .Q(U99_DATA1_6) );
  DLH_X1 round_in_key_reg_6_ ( .G(n5470), .D(U99_DATA1_6), .Q(n3398) );
  DLH_X1 expanded_key_in_reg_6_ ( .G(n5472), .D(n4451), .Q(n3139) );
  DFF_X1 expanded_key_reg_7_ ( .D(n4163), .CK(clk), .Q(U99_DATA1_7) );
  DLH_X1 round_in_key_reg_7_ ( .G(n5470), .D(U99_DATA1_7), .Q(n3399) );
  DLH_X1 expanded_key_in_reg_7_ ( .G(n5474), .D(n4450), .Q(n3140) );
  DFF_X1 expanded_key_reg_8_ ( .D(n4162), .CK(clk), .Q(U99_DATA1_8) );
  DLH_X1 round_in_key_reg_8_ ( .G(n5470), .D(U99_DATA1_8), .Q(n3400) );
  DLH_X1 expanded_key_in_reg_8_ ( .G(n5475), .D(n4449), .Q(n3141) );
  DFF_X1 expanded_key_reg_9_ ( .D(n4161), .CK(clk), .Q(U99_DATA1_9) );
  DLH_X1 round_in_key_reg_9_ ( .G(n5470), .D(U99_DATA1_9), .Q(n3401) );
  DLH_X1 expanded_key_in_reg_9_ ( .G(n5472), .D(n4448), .Q(n3142) );
  DFF_X1 expanded_key_reg_10_ ( .D(n4160), .CK(clk), .Q(U99_DATA1_10) );
  DLH_X1 round_in_key_reg_10_ ( .G(n5470), .D(U99_DATA1_10), .Q(n3402) );
  DLH_X1 expanded_key_in_reg_10_ ( .G(U47_Z_1), .D(n4447), .Q(n3143) );
  DFF_X1 expanded_key_reg_11_ ( .D(n4159), .CK(clk), .Q(U99_DATA1_11) );
  DLH_X1 round_in_key_reg_11_ ( .G(n5470), .D(U99_DATA1_11), .Q(n3403) );
  DLH_X1 expanded_key_in_reg_11_ ( .G(n5472), .D(n4446), .Q(n3144) );
  DFF_X1 expanded_key_reg_12_ ( .D(n4158), .CK(clk), .Q(U99_DATA1_12) );
  DLH_X1 round_in_key_reg_12_ ( .G(n5469), .D(U99_DATA1_12), .Q(n3404) );
  DLH_X1 expanded_key_in_reg_12_ ( .G(n5473), .D(n4445), .Q(n3145) );
  DFF_X1 expanded_key_reg_13_ ( .D(n4157), .CK(clk), .Q(U99_DATA1_13) );
  DLH_X1 round_in_key_reg_13_ ( .G(n5469), .D(U99_DATA1_13), .Q(n3405) );
  DLH_X1 expanded_key_in_reg_13_ ( .G(n5473), .D(n4444), .Q(n3146) );
  DFF_X1 expanded_key_reg_14_ ( .D(n4156), .CK(clk), .Q(U99_DATA1_14) );
  DLH_X1 round_in_key_reg_14_ ( .G(n5469), .D(U99_DATA1_14), .Q(n3406) );
  DLH_X1 expanded_key_in_reg_14_ ( .G(n5474), .D(n4443), .Q(n3147) );
  DFF_X1 expanded_key_reg_15_ ( .D(n4155), .CK(clk), .Q(U99_DATA1_15) );
  DLH_X1 round_in_key_reg_15_ ( .G(n5469), .D(U99_DATA1_15), .Q(n3407) );
  DLH_X1 expanded_key_in_reg_15_ ( .G(n5475), .D(n4442), .Q(n3148) );
  DFF_X1 expanded_key_reg_16_ ( .D(n4154), .CK(clk), .Q(U99_DATA1_16) );
  DLH_X1 round_in_key_reg_16_ ( .G(n5469), .D(U99_DATA1_16), .Q(n3408) );
  DLH_X1 expanded_key_in_reg_16_ ( .G(n5475), .D(n4441), .Q(n3149) );
  DFF_X1 expanded_key_reg_17_ ( .D(n4153), .CK(clk), .Q(U99_DATA1_17) );
  DLH_X1 round_in_key_reg_17_ ( .G(n5469), .D(U99_DATA1_17), .Q(n3409) );
  DLH_X1 expanded_key_in_reg_17_ ( .G(n5474), .D(n4440), .Q(n3150) );
  DFF_X1 expanded_key_reg_18_ ( .D(n4152), .CK(clk), .Q(U99_DATA1_18) );
  DLH_X1 round_in_key_reg_18_ ( .G(n5469), .D(U99_DATA1_18), .Q(n3410) );
  DLH_X1 expanded_key_in_reg_18_ ( .G(U47_Z_1), .D(n4439), .Q(n3151) );
  DFF_X1 expanded_key_reg_19_ ( .D(n4151), .CK(clk), .Q(U99_DATA1_19) );
  DLH_X1 round_in_key_reg_19_ ( .G(n5469), .D(U99_DATA1_19), .Q(n3411) );
  DLH_X1 expanded_key_in_reg_19_ ( .G(n5474), .D(n4438), .Q(n3152) );
  DFF_X1 expanded_key_reg_20_ ( .D(n4150), .CK(clk), .Q(U99_DATA1_20) );
  DLH_X1 round_in_key_reg_20_ ( .G(n5469), .D(U99_DATA1_20), .Q(n3412) );
  DLH_X1 expanded_key_in_reg_20_ ( .G(n5473), .D(n4437), .Q(n3153) );
  DFF_X1 expanded_key_reg_21_ ( .D(n4149), .CK(clk), .Q(U99_DATA1_21) );
  DLH_X1 round_in_key_reg_21_ ( .G(n5469), .D(U99_DATA1_21), .Q(n3413) );
  DLH_X1 expanded_key_in_reg_21_ ( .G(n5472), .D(n4436), .Q(n3154) );
  DFF_X1 expanded_key_reg_22_ ( .D(n4148), .CK(clk), .Q(U99_DATA1_22) );
  DLH_X1 round_in_key_reg_22_ ( .G(n5469), .D(U99_DATA1_22), .Q(n3414) );
  DLH_X1 expanded_key_in_reg_22_ ( .G(n5473), .D(n4435), .Q(n3155) );
  DFF_X1 expanded_key_reg_23_ ( .D(n4147), .CK(clk), .Q(U99_DATA1_23) );
  DLH_X1 round_in_key_reg_23_ ( .G(n5468), .D(U99_DATA1_23), .Q(n3415) );
  DLH_X1 expanded_key_in_reg_23_ ( .G(n5474), .D(n4434), .Q(n3156) );
  DFF_X1 expanded_key_reg_24_ ( .D(n4146), .CK(clk), .Q(U99_DATA1_24) );
  DLH_X1 round_in_key_reg_24_ ( .G(n5468), .D(U99_DATA1_24), .Q(n3416) );
  DLH_X1 expanded_key_in_reg_24_ ( .G(n5472), .D(n4433), .Q(n3157) );
  DFF_X1 expanded_key_reg_25_ ( .D(n4145), .CK(clk), .Q(U99_DATA1_25) );
  DLH_X1 round_in_key_reg_25_ ( .G(n5468), .D(U99_DATA1_25), .Q(n3417) );
  DLH_X1 expanded_key_in_reg_25_ ( .G(n5472), .D(n4432), .Q(n3158) );
  DFF_X1 expanded_key_reg_26_ ( .D(n4144), .CK(clk), .Q(U99_DATA1_26) );
  DLH_X1 round_in_key_reg_26_ ( .G(n5468), .D(U99_DATA1_26), .Q(n3418) );
  DLH_X1 expanded_key_in_reg_26_ ( .G(n5473), .D(n4431), .Q(n3159) );
  DFF_X1 expanded_key_reg_27_ ( .D(n4143), .CK(clk), .Q(U99_DATA1_27) );
  DLH_X1 round_in_key_reg_27_ ( .G(n5468), .D(U99_DATA1_27), .Q(n3419) );
  DLH_X1 expanded_key_in_reg_27_ ( .G(n5472), .D(n4430), .Q(n3160) );
  DFF_X1 expanded_key_reg_28_ ( .D(n4142), .CK(clk), .Q(U99_DATA1_28) );
  DLH_X1 round_in_key_reg_28_ ( .G(n5468), .D(U99_DATA1_28), .Q(n3420) );
  DLH_X1 expanded_key_in_reg_28_ ( .G(n5473), .D(n4429), .Q(n3161) );
  DFF_X1 expanded_key_reg_29_ ( .D(n4141), .CK(clk), .Q(U99_DATA1_29) );
  DLH_X1 round_in_key_reg_29_ ( .G(n5468), .D(U99_DATA1_29), .Q(n3421) );
  DLH_X1 expanded_key_in_reg_29_ ( .G(n5473), .D(n4428), .Q(n3162) );
  DFF_X1 expanded_key_reg_30_ ( .D(n4140), .CK(clk), .Q(U99_DATA1_30) );
  DLH_X1 round_in_key_reg_30_ ( .G(n5468), .D(U99_DATA1_30), .Q(n3422) );
  DLH_X1 expanded_key_in_reg_30_ ( .G(U47_Z_1), .D(n4427), .Q(n3163) );
  DFF_X1 expanded_key_reg_31_ ( .D(n4139), .CK(clk), .Q(U99_DATA1_31) );
  DLH_X1 round_in_key_reg_31_ ( .G(n5468), .D(U99_DATA1_31), .Q(n3423) );
  DLH_X1 expanded_key_in_reg_31_ ( .G(n5475), .D(n4426), .Q(n3164) );
  DFF_X1 expanded_key_reg_32_ ( .D(n4138), .CK(clk), .Q(U99_DATA1_32) );
  DLH_X1 round_in_key_reg_32_ ( .G(n5468), .D(U99_DATA1_32), .Q(n3424) );
  DLH_X1 expanded_key_in_reg_32_ ( .G(n5475), .D(n4425), .Q(n3165) );
  DFF_X1 expanded_key_reg_33_ ( .D(n4137), .CK(clk), .Q(U99_DATA1_33) );
  DLH_X1 round_in_key_reg_33_ ( .G(n5468), .D(U99_DATA1_33), .Q(n3425) );
  DLH_X1 expanded_key_in_reg_33_ ( .G(n5473), .D(n4424), .Q(n3166) );
  DFF_X1 expanded_key_reg_34_ ( .D(n4136), .CK(clk), .Q(U99_DATA1_34) );
  DLH_X1 round_in_key_reg_34_ ( .G(n5467), .D(U99_DATA1_34), .Q(n3426) );
  DLH_X1 expanded_key_in_reg_34_ ( .G(n5475), .D(n4423), .Q(n3167) );
  DFF_X1 expanded_key_reg_35_ ( .D(n4135), .CK(clk), .Q(U99_DATA1_35) );
  DLH_X1 round_in_key_reg_35_ ( .G(n5467), .D(U99_DATA1_35), .Q(n3427) );
  DLH_X1 expanded_key_in_reg_35_ ( .G(n5472), .D(n4422), .Q(n3168) );
  DFF_X1 expanded_key_reg_36_ ( .D(n4134), .CK(clk), .Q(U99_DATA1_36) );
  DLH_X1 round_in_key_reg_36_ ( .G(n5467), .D(U99_DATA1_36), .Q(n3428) );
  DLH_X1 expanded_key_in_reg_36_ ( .G(n5472), .D(n4421), .Q(n3169) );
  DFF_X1 expanded_key_reg_37_ ( .D(n4133), .CK(clk), .Q(U99_DATA1_37) );
  DLH_X1 round_in_key_reg_37_ ( .G(n5467), .D(U99_DATA1_37), .Q(n3429) );
  DLH_X1 expanded_key_in_reg_37_ ( .G(n5474), .D(n4420), .Q(n3170) );
  DFF_X1 expanded_key_reg_38_ ( .D(n4132), .CK(clk), .Q(U99_DATA1_38) );
  DLH_X1 round_in_key_reg_38_ ( .G(n5467), .D(U99_DATA1_38), .Q(n3430) );
  DLH_X1 expanded_key_in_reg_38_ ( .G(n5472), .D(n4419), .Q(n3171) );
  DFF_X1 expanded_key_reg_39_ ( .D(n4131), .CK(clk), .Q(U99_DATA1_39) );
  DLH_X1 round_in_key_reg_39_ ( .G(n5467), .D(U99_DATA1_39), .Q(n3431) );
  DLH_X1 expanded_key_in_reg_39_ ( .G(n5475), .D(n4418), .Q(n3172) );
  DFF_X1 expanded_key_reg_40_ ( .D(n4130), .CK(clk), .Q(U99_DATA1_40) );
  DLH_X1 round_in_key_reg_40_ ( .G(n5467), .D(U99_DATA1_40), .Q(n3432) );
  DLH_X1 expanded_key_in_reg_40_ ( .G(n5475), .D(n4417), .Q(n3173) );
  DFF_X1 expanded_key_reg_41_ ( .D(n4129), .CK(clk), .Q(U99_DATA1_41) );
  DLH_X1 round_in_key_reg_41_ ( .G(n5467), .D(U99_DATA1_41), .Q(n3433) );
  DLH_X1 expanded_key_in_reg_41_ ( .G(n5475), .D(n4416), .Q(n3174) );
  DFF_X1 expanded_key_reg_42_ ( .D(n4128), .CK(clk), .Q(U99_DATA1_42) );
  DLH_X1 round_in_key_reg_42_ ( .G(n5467), .D(U99_DATA1_42), .Q(n3434) );
  DLH_X1 expanded_key_in_reg_42_ ( .G(n5475), .D(n4415), .Q(n3175) );
  DFF_X1 expanded_key_reg_43_ ( .D(n4127), .CK(clk), .Q(U99_DATA1_43) );
  DLH_X1 round_in_key_reg_43_ ( .G(n5467), .D(U99_DATA1_43), .Q(n3435) );
  DLH_X1 expanded_key_in_reg_43_ ( .G(n5475), .D(n4414), .Q(n3176) );
  DFF_X1 expanded_key_reg_44_ ( .D(n4126), .CK(clk), .Q(U99_DATA1_44) );
  DLH_X1 round_in_key_reg_44_ ( .G(n5467), .D(U99_DATA1_44), .Q(n3436) );
  DLH_X1 expanded_key_in_reg_44_ ( .G(n5475), .D(n4413), .Q(n3177) );
  DFF_X1 expanded_key_reg_45_ ( .D(n4125), .CK(clk), .Q(U99_DATA1_45) );
  DLH_X1 round_in_key_reg_45_ ( .G(n5466), .D(U99_DATA1_45), .Q(n3437) );
  DLH_X1 expanded_key_in_reg_45_ ( .G(n5475), .D(n4412), .Q(n3178) );
  DFF_X1 expanded_key_reg_46_ ( .D(n4124), .CK(clk), .Q(U99_DATA1_46) );
  DLH_X1 round_in_key_reg_46_ ( .G(n5466), .D(U99_DATA1_46), .Q(n3438) );
  DLH_X1 expanded_key_in_reg_46_ ( .G(n5475), .D(n4411), .Q(n3179) );
  DFF_X1 expanded_key_reg_47_ ( .D(n4123), .CK(clk), .Q(U99_DATA1_47) );
  DLH_X1 round_in_key_reg_47_ ( .G(n5466), .D(U99_DATA1_47), .Q(n3439) );
  DLH_X1 expanded_key_in_reg_47_ ( .G(n5475), .D(n4410), .Q(n3180) );
  DFF_X1 expanded_key_reg_48_ ( .D(n4122), .CK(clk), .Q(U99_DATA1_48) );
  DLH_X1 round_in_key_reg_48_ ( .G(n5466), .D(U99_DATA1_48), .Q(n3440) );
  DLH_X1 expanded_key_in_reg_48_ ( .G(n5475), .D(n4409), .Q(n3181) );
  DFF_X1 expanded_key_reg_49_ ( .D(n4121), .CK(clk), .Q(U99_DATA1_49) );
  DLH_X1 round_in_key_reg_49_ ( .G(n5466), .D(U99_DATA1_49), .Q(n3441) );
  DLH_X1 expanded_key_in_reg_49_ ( .G(n5475), .D(n4408), .Q(n3182) );
  DFF_X1 expanded_key_reg_50_ ( .D(n4120), .CK(clk), .Q(U99_DATA1_50) );
  DLH_X1 round_in_key_reg_50_ ( .G(n5466), .D(U99_DATA1_50), .Q(n3442) );
  DLH_X1 expanded_key_in_reg_50_ ( .G(n5474), .D(n4407), .Q(n3183) );
  DFF_X1 expanded_key_reg_51_ ( .D(n4119), .CK(clk), .Q(U99_DATA1_51) );
  DLH_X1 round_in_key_reg_51_ ( .G(n5466), .D(U99_DATA1_51), .Q(n3443) );
  DLH_X1 expanded_key_in_reg_51_ ( .G(n5474), .D(n4406), .Q(n3184) );
  DFF_X1 expanded_key_reg_52_ ( .D(n4118), .CK(clk), .Q(U99_DATA1_52) );
  DLH_X1 round_in_key_reg_52_ ( .G(n5466), .D(U99_DATA1_52), .Q(n3444) );
  DLH_X1 expanded_key_in_reg_52_ ( .G(n5474), .D(n4405), .Q(n3185) );
  DFF_X1 expanded_key_reg_53_ ( .D(n4117), .CK(clk), .Q(U99_DATA1_53) );
  DLH_X1 round_in_key_reg_53_ ( .G(n5466), .D(U99_DATA1_53), .Q(n3445) );
  DLH_X1 expanded_key_in_reg_53_ ( .G(n5474), .D(n4404), .Q(n3186) );
  DFF_X1 expanded_key_reg_54_ ( .D(n4116), .CK(clk), .Q(U99_DATA1_54) );
  DLH_X1 round_in_key_reg_54_ ( .G(n5466), .D(U99_DATA1_54), .Q(n3446) );
  DLH_X1 expanded_key_in_reg_54_ ( .G(n5474), .D(n4403), .Q(n3187) );
  DFF_X1 expanded_key_reg_55_ ( .D(n4115), .CK(clk), .Q(U99_DATA1_55) );
  DLH_X1 round_in_key_reg_55_ ( .G(n5466), .D(U99_DATA1_55), .Q(n3447) );
  DLH_X1 expanded_key_in_reg_55_ ( .G(n5474), .D(n4402), .Q(n3188) );
  DFF_X1 expanded_key_reg_56_ ( .D(n4114), .CK(clk), .Q(U99_DATA1_56) );
  DLH_X1 round_in_key_reg_56_ ( .G(n5468), .D(U99_DATA1_56), .Q(n3448) );
  DLH_X1 expanded_key_in_reg_56_ ( .G(n5474), .D(n4401), .Q(n3189) );
  DFF_X1 expanded_key_reg_57_ ( .D(n4113), .CK(clk), .Q(U99_DATA1_57) );
  DLH_X1 round_in_key_reg_57_ ( .G(n5468), .D(U99_DATA1_57), .Q(n3449) );
  DLH_X1 expanded_key_in_reg_57_ ( .G(n5474), .D(n4400), .Q(n3190) );
  DFF_X1 expanded_key_reg_58_ ( .D(n4112), .CK(clk), .Q(U99_DATA1_58) );
  DLH_X1 round_in_key_reg_58_ ( .G(n5466), .D(U99_DATA1_58), .Q(n3450) );
  DLH_X1 expanded_key_in_reg_58_ ( .G(n5474), .D(n4399), .Q(n3191) );
  DFF_X1 expanded_key_reg_59_ ( .D(n4111), .CK(clk), .Q(U99_DATA1_59) );
  DLH_X1 round_in_key_reg_59_ ( .G(n5471), .D(U99_DATA1_59), .Q(n3451) );
  DLH_X1 expanded_key_in_reg_59_ ( .G(n5474), .D(n4398), .Q(n3192) );
  DFF_X1 expanded_key_reg_60_ ( .D(n4110), .CK(clk), .Q(U99_DATA1_60) );
  DLH_X1 round_in_key_reg_60_ ( .G(n5464), .D(U99_DATA1_60), .Q(n3452) );
  DLH_X1 expanded_key_in_reg_60_ ( .G(n5474), .D(n4397), .Q(n3193) );
  DFF_X1 expanded_key_reg_61_ ( .D(n4109), .CK(clk), .Q(U99_DATA1_61) );
  DLH_X1 round_in_key_reg_61_ ( .G(n5470), .D(U99_DATA1_61), .Q(n3453) );
  DLH_X1 expanded_key_in_reg_61_ ( .G(n5473), .D(n4396), .Q(n3194) );
  DFF_X1 expanded_key_reg_62_ ( .D(n4108), .CK(clk), .Q(U99_DATA1_62) );
  DLH_X1 round_in_key_reg_62_ ( .G(n5470), .D(U99_DATA1_62), .Q(n3454) );
  DLH_X1 expanded_key_in_reg_62_ ( .G(U47_Z_1), .D(n4395), .Q(n3195) );
  DFF_X1 expanded_key_reg_63_ ( .D(n4107), .CK(clk), .Q(U99_DATA1_63) );
  DLH_X1 round_in_key_reg_63_ ( .G(n5465), .D(U99_DATA1_63), .Q(n3455) );
  DLH_X1 expanded_key_in_reg_63_ ( .G(U47_Z_1), .D(n4394), .Q(n3196) );
  DFF_X1 expanded_key_reg_64_ ( .D(n4106), .CK(clk), .Q(U99_DATA1_64) );
  DLH_X1 round_in_key_reg_64_ ( .G(n5468), .D(U99_DATA1_64), .Q(n3456) );
  DLH_X1 expanded_key_in_reg_64_ ( .G(n5473), .D(n4393), .Q(n3197) );
  DFF_X1 expanded_key_reg_65_ ( .D(n4105), .CK(clk), .Q(U99_DATA1_65) );
  DLH_X1 round_in_key_reg_65_ ( .G(n5469), .D(U99_DATA1_65), .Q(n3457) );
  DLH_X1 expanded_key_in_reg_65_ ( .G(U47_Z_1), .D(n4392), .Q(n3198) );
  DFF_X1 expanded_key_reg_66_ ( .D(n4104), .CK(clk), .Q(U99_DATA1_66) );
  DLH_X1 round_in_key_reg_66_ ( .G(n5467), .D(U99_DATA1_66), .Q(n3458) );
  DLH_X1 expanded_key_in_reg_66_ ( .G(U47_Z_1), .D(n4391), .Q(n3199) );
  DFF_X1 expanded_key_reg_67_ ( .D(n4103), .CK(clk), .Q(U99_DATA1_67) );
  DLH_X1 round_in_key_reg_67_ ( .G(n5465), .D(U99_DATA1_67), .Q(n3459) );
  DLH_X1 expanded_key_in_reg_67_ ( .G(U47_Z_1), .D(n4390), .Q(n3200) );
  DFF_X1 expanded_key_reg_68_ ( .D(n4102), .CK(clk), .Q(U99_DATA1_68) );
  DLH_X1 round_in_key_reg_68_ ( .G(n5471), .D(U99_DATA1_68), .Q(n3460) );
  DLH_X1 expanded_key_in_reg_68_ ( .G(U47_Z_1), .D(n4389), .Q(n3201) );
  DFF_X1 expanded_key_reg_69_ ( .D(n4101), .CK(clk), .Q(U99_DATA1_69) );
  DLH_X1 round_in_key_reg_69_ ( .G(n5470), .D(U99_DATA1_69), .Q(n3461) );
  DLH_X1 expanded_key_in_reg_69_ ( .G(n5472), .D(n4388), .Q(n3202) );
  DFF_X1 expanded_key_reg_70_ ( .D(n4100), .CK(clk), .Q(U99_DATA1_70) );
  DLH_X1 round_in_key_reg_70_ ( .G(n5466), .D(U99_DATA1_70), .Q(n3462) );
  DLH_X1 expanded_key_in_reg_70_ ( .G(U47_Z_1), .D(n4387), .Q(n3203) );
  DFF_X1 expanded_key_reg_71_ ( .D(n4099), .CK(clk), .Q(U99_DATA1_71) );
  DLH_X1 round_in_key_reg_71_ ( .G(n5468), .D(U99_DATA1_71), .Q(n3463) );
  DLH_X1 expanded_key_in_reg_71_ ( .G(n5475), .D(n4386), .Q(n3204) );
  DFF_X1 expanded_key_reg_72_ ( .D(n4098), .CK(clk), .Q(U99_DATA1_72) );
  DLH_X1 round_in_key_reg_72_ ( .G(n5469), .D(U99_DATA1_72), .Q(n3464) );
  DLH_X1 expanded_key_in_reg_72_ ( .G(n5473), .D(n4385), .Q(n3205) );
  DFF_X1 expanded_key_reg_73_ ( .D(n4097), .CK(clk), .Q(U99_DATA1_73) );
  DLH_X1 round_in_key_reg_73_ ( .G(n5464), .D(U99_DATA1_73), .Q(n3465) );
  DLH_X1 expanded_key_in_reg_73_ ( .G(n5473), .D(n4384), .Q(n3206) );
  DFF_X1 expanded_key_reg_74_ ( .D(n4096), .CK(clk), .Q(U99_DATA1_74) );
  DLH_X1 round_in_key_reg_74_ ( .G(n5469), .D(U99_DATA1_74), .Q(n3466) );
  DLH_X1 expanded_key_in_reg_74_ ( .G(n5473), .D(n4383), .Q(n3207) );
  DFF_X1 expanded_key_reg_75_ ( .D(n4095), .CK(clk), .Q(U99_DATA1_75) );
  DLH_X1 round_in_key_reg_75_ ( .G(n5470), .D(U99_DATA1_75), .Q(n3467) );
  DLH_X1 expanded_key_in_reg_75_ ( .G(n5473), .D(n4382), .Q(n3208) );
  DFF_X1 expanded_key_reg_76_ ( .D(n4094), .CK(clk), .Q(U99_DATA1_76) );
  DLH_X1 round_in_key_reg_76_ ( .G(n5467), .D(U99_DATA1_76), .Q(n3468) );
  DLH_X1 expanded_key_in_reg_76_ ( .G(n5473), .D(n4381), .Q(n3209) );
  DFF_X1 expanded_key_reg_77_ ( .D(n4093), .CK(clk), .Q(U99_DATA1_77) );
  DLH_X1 round_in_key_reg_77_ ( .G(n5467), .D(U99_DATA1_77), .Q(n3469) );
  DLH_X1 expanded_key_in_reg_77_ ( .G(n5473), .D(n4380), .Q(n3210) );
  DFF_X1 expanded_key_reg_78_ ( .D(n4092), .CK(clk), .Q(U99_DATA1_78) );
  DLH_X1 round_in_key_reg_78_ ( .G(n5466), .D(U99_DATA1_78), .Q(n3470) );
  DLH_X1 expanded_key_in_reg_78_ ( .G(n5473), .D(n4379), .Q(n3211) );
  DFF_X1 expanded_key_reg_79_ ( .D(n4091), .CK(clk), .Q(U99_DATA1_79) );
  DLH_X1 round_in_key_reg_79_ ( .G(n5464), .D(U99_DATA1_79), .Q(n3471) );
  DLH_X1 expanded_key_in_reg_79_ ( .G(n5473), .D(n4378), .Q(n3212) );
  DFF_X1 expanded_key_reg_80_ ( .D(n4090), .CK(clk), .Q(U99_DATA1_80) );
  DLH_X1 round_in_key_reg_80_ ( .G(n5467), .D(U99_DATA1_80), .Q(n3472) );
  DLH_X1 expanded_key_in_reg_80_ ( .G(n5473), .D(n4377), .Q(n3213) );
  DFF_X1 expanded_key_reg_81_ ( .D(n4089), .CK(clk), .Q(U99_DATA1_81) );
  DLH_X1 round_in_key_reg_81_ ( .G(n5468), .D(U99_DATA1_81), .Q(n3473) );
  DLH_X1 expanded_key_in_reg_81_ ( .G(n5473), .D(n4376), .Q(n3214) );
  DFF_X1 expanded_key_reg_82_ ( .D(n4088), .CK(clk), .Q(U99_DATA1_82) );
  DLH_X1 round_in_key_reg_82_ ( .G(n5465), .D(U99_DATA1_82), .Q(n3474) );
  DLH_X1 expanded_key_in_reg_82_ ( .G(n5473), .D(n4375), .Q(n3215) );
  DFF_X1 expanded_key_reg_83_ ( .D(n4087), .CK(clk), .Q(U99_DATA1_83) );
  DLH_X1 round_in_key_reg_83_ ( .G(n5468), .D(U99_DATA1_83), .Q(n3475) );
  DLH_X1 expanded_key_in_reg_83_ ( .G(n5472), .D(n4374), .Q(n3216) );
  DFF_X1 expanded_key_reg_84_ ( .D(n4086), .CK(clk), .Q(U99_DATA1_84) );
  DLH_X1 round_in_key_reg_84_ ( .G(n5470), .D(U99_DATA1_84), .Q(n3476) );
  DLH_X1 expanded_key_in_reg_84_ ( .G(n5472), .D(n4373), .Q(n3217) );
  DFF_X1 expanded_key_reg_85_ ( .D(n4085), .CK(clk), .Q(U99_DATA1_85) );
  DLH_X1 round_in_key_reg_85_ ( .G(n5469), .D(U99_DATA1_85), .Q(n3477) );
  DLH_X1 expanded_key_in_reg_85_ ( .G(n5472), .D(n4372), .Q(n3218) );
  DFF_X1 expanded_key_reg_86_ ( .D(n4084), .CK(clk), .Q(U99_DATA1_86) );
  DLH_X1 round_in_key_reg_86_ ( .G(n5469), .D(U99_DATA1_86), .Q(n3478) );
  DLH_X1 expanded_key_in_reg_86_ ( .G(n5472), .D(n4371), .Q(n3219) );
  DFF_X1 expanded_key_reg_87_ ( .D(n4083), .CK(clk), .Q(U99_DATA1_87) );
  DLH_X1 round_in_key_reg_87_ ( .G(n5468), .D(U99_DATA1_87), .Q(n3479) );
  DLH_X1 expanded_key_in_reg_87_ ( .G(n5472), .D(n4370), .Q(n3220) );
  DFF_X1 expanded_key_reg_88_ ( .D(n4082), .CK(clk), .Q(U99_DATA1_88) );
  DLH_X1 round_in_key_reg_88_ ( .G(n5466), .D(U99_DATA1_88), .Q(n3480) );
  DLH_X1 expanded_key_in_reg_88_ ( .G(n5472), .D(n4369), .Q(n3221) );
  DFF_X1 expanded_key_reg_89_ ( .D(n4081), .CK(clk), .Q(U99_DATA1_89) );
  DLH_X1 round_in_key_reg_89_ ( .G(n5464), .D(U99_DATA1_89), .Q(n3481) );
  DLH_X1 expanded_key_in_reg_89_ ( .G(n5472), .D(n4368), .Q(n3222) );
  DFF_X1 expanded_key_reg_90_ ( .D(n4080), .CK(clk), .Q(U99_DATA1_90) );
  DLH_X1 round_in_key_reg_90_ ( .G(n5465), .D(U99_DATA1_90), .Q(n3482) );
  DLH_X1 expanded_key_in_reg_90_ ( .G(n5472), .D(n4367), .Q(n3223) );
  DFF_X1 expanded_key_reg_91_ ( .D(n4079), .CK(clk), .Q(U99_DATA1_91) );
  DLH_X1 round_in_key_reg_91_ ( .G(n5467), .D(U99_DATA1_91), .Q(n3483) );
  DLH_X1 expanded_key_in_reg_91_ ( .G(n5472), .D(n4366), .Q(n3224) );
  DFF_X1 expanded_key_reg_92_ ( .D(n4078), .CK(clk), .Q(U99_DATA1_92) );
  DLH_X1 round_in_key_reg_92_ ( .G(n5470), .D(U99_DATA1_92), .Q(n3484) );
  DLH_X1 expanded_key_in_reg_92_ ( .G(n5472), .D(n4365), .Q(n3225) );
  DFF_X1 expanded_key_reg_93_ ( .D(n4077), .CK(clk), .Q(U99_DATA1_93) );
  DLH_X1 round_in_key_reg_93_ ( .G(n5469), .D(U99_DATA1_93), .Q(n3485) );
  DLH_X1 expanded_key_in_reg_93_ ( .G(n5472), .D(n4364), .Q(n3226) );
  DFF_X1 expanded_key_reg_94_ ( .D(n4076), .CK(clk), .Q(U99_DATA1_94) );
  DLH_X1 round_in_key_reg_94_ ( .G(n5464), .D(U99_DATA1_94), .Q(n3486) );
  DLH_X1 expanded_key_in_reg_94_ ( .G(n5475), .D(n4363), .Q(n3227) );
  DFF_X1 expanded_key_reg_95_ ( .D(n4075), .CK(clk), .Q(U99_DATA1_95) );
  DLH_X1 round_in_key_reg_95_ ( .G(n5464), .D(U99_DATA1_95), .Q(n3487) );
  DLH_X1 expanded_key_in_reg_95_ ( .G(n5475), .D(n4362), .Q(n3228) );
  DFF_X1 expanded_key_reg_96_ ( .D(n4074), .CK(clk), .Q(U99_DATA1_96) );
  DLH_X1 round_in_key_reg_96_ ( .G(n5466), .D(U99_DATA1_96), .Q(n3488) );
  DLH_X1 expanded_key_in_reg_96_ ( .G(n5473), .D(n4361), .Q(n3229) );
  DFF_X1 expanded_key_reg_97_ ( .D(n4073), .CK(clk), .Q(U99_DATA1_97) );
  DLH_X1 round_in_key_reg_97_ ( .G(n5467), .D(U99_DATA1_97), .Q(n3489) );
  DLH_X1 expanded_key_in_reg_97_ ( .G(n5474), .D(n4360), .Q(n3230) );
  DFF_X1 expanded_key_reg_98_ ( .D(n4072), .CK(clk), .Q(U99_DATA1_98) );
  DLH_X1 round_in_key_reg_98_ ( .G(n5471), .D(U99_DATA1_98), .Q(n3490) );
  DLH_X1 expanded_key_in_reg_98_ ( .G(n5472), .D(n4359), .Q(n3231) );
  DFF_X1 expanded_key_reg_99_ ( .D(n4198), .CK(clk), .Q(U99_DATA1_99) );
  DLH_X1 round_in_key_reg_99_ ( .G(n5468), .D(U99_DATA1_99), .Q(n3491) );
  DLH_X1 expanded_key_in_reg_99_ ( .G(n5472), .D(n4358), .Q(n3232) );
  DFF_X1 expanded_key_reg_100_ ( .D(n4197), .CK(clk), .Q(U99_DATA1_100) );
  DLH_X1 round_in_key_reg_100_ ( .G(n5470), .D(U99_DATA1_100), .Q(n3492) );
  DLH_X1 expanded_key_in_reg_100_ ( .G(n5473), .D(n4357), .Q(n3233) );
  DFF_X1 expanded_key_reg_101_ ( .D(n4196), .CK(clk), .Q(U99_DATA1_101) );
  DLH_X1 round_in_key_reg_101_ ( .G(n5467), .D(U99_DATA1_101), .Q(n3493) );
  DLH_X1 expanded_key_in_reg_101_ ( .G(U47_Z_1), .D(n4356), .Q(n3234) );
  DFF_X1 expanded_key_reg_102_ ( .D(n4195), .CK(clk), .Q(U99_DATA1_102) );
  DLH_X1 round_in_key_reg_102_ ( .G(n5465), .D(U99_DATA1_102), .Q(n3494) );
  DLH_X1 expanded_key_in_reg_102_ ( .G(U47_Z_1), .D(n4355), .Q(n3235) );
  DFF_X1 expanded_key_reg_103_ ( .D(n4194), .CK(clk), .Q(U99_DATA1_103) );
  DLH_X1 round_in_key_reg_103_ ( .G(n5464), .D(U99_DATA1_103), .Q(n3495) );
  DLH_X1 expanded_key_in_reg_103_ ( .G(n5474), .D(n4354), .Q(n3236) );
  DFF_X1 expanded_key_reg_104_ ( .D(n4193), .CK(clk), .Q(U99_DATA1_104) );
  DLH_X1 round_in_key_reg_104_ ( .G(n5464), .D(U99_DATA1_104), .Q(n3496) );
  DLH_X1 expanded_key_in_reg_104_ ( .G(n5475), .D(n4353), .Q(n3237) );
  DFF_X1 expanded_key_reg_105_ ( .D(n4192), .CK(clk), .Q(U99_DATA1_105) );
  DLH_X1 round_in_key_reg_105_ ( .G(n5466), .D(U99_DATA1_105), .Q(n3497) );
  DLH_X1 expanded_key_in_reg_105_ ( .G(n5475), .D(n4352), .Q(n3238) );
  DFF_X1 expanded_key_reg_106_ ( .D(n4191), .CK(clk), .Q(U99_DATA1_106) );
  DLH_X1 round_in_key_reg_106_ ( .G(n5465), .D(U99_DATA1_106), .Q(n3498) );
  DLH_X1 expanded_key_in_reg_106_ ( .G(n5475), .D(n4351), .Q(n3239) );
  DFF_X1 expanded_key_reg_107_ ( .D(n4190), .CK(clk), .Q(U99_DATA1_107) );
  DLH_X1 round_in_key_reg_107_ ( .G(n5466), .D(U99_DATA1_107), .Q(n3499) );
  DLH_X1 expanded_key_in_reg_107_ ( .G(n5475), .D(n4350), .Q(n3240) );
  DFF_X1 expanded_key_reg_108_ ( .D(n4189), .CK(clk), .Q(U99_DATA1_108) );
  DLH_X1 round_in_key_reg_108_ ( .G(n5469), .D(U99_DATA1_108), .Q(n3500) );
  DLH_X1 expanded_key_in_reg_108_ ( .G(n5475), .D(n4349), .Q(n3241) );
  DFF_X1 expanded_key_reg_109_ ( .D(n4188), .CK(clk), .Q(U99_DATA1_109) );
  DLH_X1 round_in_key_reg_109_ ( .G(n5468), .D(U99_DATA1_109), .Q(n3501) );
  DLH_X1 expanded_key_in_reg_109_ ( .G(n5474), .D(n4348), .Q(n3242) );
  DFF_X1 expanded_key_reg_110_ ( .D(n4187), .CK(clk), .Q(U99_DATA1_110) );
  DLH_X1 round_in_key_reg_110_ ( .G(n5467), .D(U99_DATA1_110), .Q(n3502) );
  DLH_X1 expanded_key_in_reg_110_ ( .G(n5474), .D(n4347), .Q(n3243) );
  DFF_X1 expanded_key_reg_111_ ( .D(n4186), .CK(clk), .Q(U99_DATA1_111) );
  DLH_X1 round_in_key_reg_111_ ( .G(n5465), .D(U99_DATA1_111), .Q(n3503) );
  DLH_X1 expanded_key_in_reg_111_ ( .G(n5474), .D(n4346), .Q(n3244) );
  DFF_X1 expanded_key_reg_112_ ( .D(n4185), .CK(clk), .Q(U99_DATA1_112) );
  DLH_X1 round_in_key_reg_112_ ( .G(n5465), .D(U99_DATA1_112), .Q(n3504) );
  DLH_X1 expanded_key_in_reg_112_ ( .G(n5475), .D(n4345), .Q(n3245) );
  DFF_X1 expanded_key_reg_113_ ( .D(n4184), .CK(clk), .Q(U99_DATA1_113) );
  DLH_X1 round_in_key_reg_113_ ( .G(n5465), .D(U99_DATA1_113), .Q(n3505) );
  DLH_X1 expanded_key_in_reg_113_ ( .G(n5474), .D(n4344), .Q(n3246) );
  DFF_X1 expanded_key_reg_114_ ( .D(n4183), .CK(clk), .Q(U99_DATA1_114) );
  DLH_X1 round_in_key_reg_114_ ( .G(n5465), .D(U99_DATA1_114), .Q(n3506) );
  DLH_X1 expanded_key_in_reg_114_ ( .G(n5474), .D(n4343), .Q(n3247) );
  DFF_X1 expanded_key_reg_115_ ( .D(n4182), .CK(clk), .Q(U99_DATA1_115) );
  DLH_X1 round_in_key_reg_115_ ( .G(n5465), .D(U99_DATA1_115), .Q(n3507) );
  DLH_X1 expanded_key_in_reg_115_ ( .G(n5474), .D(n4342), .Q(n3248) );
  DFF_X1 expanded_key_reg_116_ ( .D(n4181), .CK(clk), .Q(U99_DATA1_116) );
  DLH_X1 round_in_key_reg_116_ ( .G(n5465), .D(U99_DATA1_116), .Q(n3508) );
  DLH_X1 expanded_key_in_reg_116_ ( .G(n5473), .D(n4341), .Q(n3249) );
  DFF_X1 expanded_key_reg_117_ ( .D(n4180), .CK(clk), .Q(U99_DATA1_117) );
  DLH_X1 round_in_key_reg_117_ ( .G(n5465), .D(U99_DATA1_117), .Q(n3509) );
  DLH_X1 expanded_key_in_reg_117_ ( .G(n5472), .D(n4340), .Q(n3250) );
  DFF_X1 expanded_key_reg_118_ ( .D(n4179), .CK(clk), .Q(U99_DATA1_118) );
  DLH_X1 round_in_key_reg_118_ ( .G(n5465), .D(U99_DATA1_118), .Q(n3510) );
  DLH_X1 expanded_key_in_reg_118_ ( .G(n5475), .D(n4339), .Q(n3251) );
  DFF_X1 expanded_key_reg_119_ ( .D(n4178), .CK(clk), .Q(U99_DATA1_119) );
  DLH_X1 round_in_key_reg_119_ ( .G(n5465), .D(U99_DATA1_119), .Q(n3511) );
  DLH_X1 expanded_key_in_reg_119_ ( .G(n5473), .D(n4338), .Q(n3252) );
  DFF_X1 expanded_key_reg_120_ ( .D(n4177), .CK(clk), .Q(U99_DATA1_120) );
  DLH_X1 round_in_key_reg_120_ ( .G(n5465), .D(U99_DATA1_120), .Q(n3512) );
  DLH_X1 expanded_key_in_reg_120_ ( .G(n5473), .D(n4337), .Q(n3253) );
  DFF_X1 expanded_key_reg_121_ ( .D(n4176), .CK(clk), .Q(U99_DATA1_121) );
  DLH_X1 round_in_key_reg_121_ ( .G(n5465), .D(U99_DATA1_121), .Q(n3513) );
  DLH_X1 expanded_key_in_reg_121_ ( .G(n5474), .D(n4336), .Q(n3254) );
  DFF_X1 expanded_key_reg_122_ ( .D(n4175), .CK(clk), .Q(U99_DATA1_122) );
  DLH_X1 round_in_key_reg_122_ ( .G(n5465), .D(U99_DATA1_122), .Q(n3514) );
  DLH_X1 expanded_key_in_reg_122_ ( .G(n5472), .D(n4335), .Q(n3255) );
  DFF_X1 expanded_key_reg_123_ ( .D(n4174), .CK(clk), .Q(U99_DATA1_123) );
  DLH_X1 round_in_key_reg_123_ ( .G(n5471), .D(U99_DATA1_123), .Q(n3515) );
  DLH_X1 expanded_key_in_reg_123_ ( .G(n5474), .D(n4334), .Q(n3256) );
  DFF_X1 expanded_key_reg_124_ ( .D(n4173), .CK(clk), .Q(U99_DATA1_124) );
  DLH_X1 round_in_key_reg_124_ ( .G(n5464), .D(U99_DATA1_124), .Q(n3516) );
  DLH_X1 expanded_key_in_reg_124_ ( .G(n5475), .D(n4333), .Q(n3257) );
  DFF_X1 expanded_key_reg_125_ ( .D(n4172), .CK(clk), .Q(U99_DATA1_125) );
  DLH_X1 round_in_key_reg_125_ ( .G(n5464), .D(U99_DATA1_125), .Q(n3517) );
  DLH_X1 expanded_key_in_reg_125_ ( .G(n5475), .D(n4332), .Q(n3258) );
  DFF_X1 expanded_key_reg_126_ ( .D(n4171), .CK(clk), .Q(U99_DATA1_126) );
  DLH_X1 round_in_key_reg_126_ ( .G(n5471), .D(U99_DATA1_126), .Q(n3518) );
  DLH_X1 expanded_key_in_reg_126_ ( .G(n5474), .D(n4331), .Q(n3259) );
  DFF_X1 temp_round_data_reg_0_ ( .D(n5400), .CK(clk), .QN(n4589) );
  DLH_X1 round_in_data_reg_0_ ( .G(U46_Z_1), .D(U49_Z_0), .Q(n3520) );
  DFF_X1 cipher_text_reg_0_ ( .D(n5401), .CK(clk), .Q(out_data[0]) );
  DFF_X1 temp_round_data_reg_1_ ( .D(n5398), .CK(clk), .QN(n4588) );
  DLH_X1 round_in_data_reg_1_ ( .G(n5471), .D(U49_Z_1), .Q(n3521) );
  DFF_X1 cipher_text_reg_1_ ( .D(n5399), .CK(clk), .Q(out_data[1]) );
  DFF_X1 temp_round_data_reg_2_ ( .D(n5396), .CK(clk), .QN(n4587) );
  DLH_X1 round_in_data_reg_2_ ( .G(U46_Z_1), .D(U49_Z_2), .Q(n3522) );
  DFF_X1 cipher_text_reg_2_ ( .D(n5397), .CK(clk), .Q(out_data[2]) );
  DFF_X1 temp_round_data_reg_3_ ( .D(n5394), .CK(clk), .QN(n4586) );
  DLH_X1 round_in_data_reg_3_ ( .G(n5466), .D(U49_Z_3), .Q(n3523) );
  DFF_X1 cipher_text_reg_3_ ( .D(n5395), .CK(clk), .Q(out_data[3]) );
  DFF_X1 temp_round_data_reg_4_ ( .D(n5392), .CK(clk), .QN(n4585) );
  DLH_X1 round_in_data_reg_4_ ( .G(n5464), .D(U49_Z_4), .Q(n3524) );
  DFF_X1 cipher_text_reg_4_ ( .D(n5393), .CK(clk), .Q(out_data[4]) );
  DFF_X1 temp_round_data_reg_5_ ( .D(n5390), .CK(clk), .QN(n4584) );
  DLH_X1 round_in_data_reg_5_ ( .G(n5467), .D(U49_Z_5), .Q(n3525) );
  DFF_X1 cipher_text_reg_5_ ( .D(n5391), .CK(clk), .Q(out_data[5]) );
  DFF_X1 temp_round_data_reg_6_ ( .D(n5388), .CK(clk), .QN(n4583) );
  DLH_X1 round_in_data_reg_6_ ( .G(n5464), .D(U49_Z_6), .Q(n3526) );
  DFF_X1 cipher_text_reg_6_ ( .D(n5389), .CK(clk), .Q(out_data[6]) );
  DFF_X1 temp_round_data_reg_7_ ( .D(n5386), .CK(clk), .QN(n4582) );
  DLH_X1 round_in_data_reg_7_ ( .G(U46_Z_1), .D(U49_Z_7), .Q(n3527) );
  DFF_X1 cipher_text_reg_7_ ( .D(n5387), .CK(clk), .Q(out_data[7]) );
  DFF_X1 temp_round_data_reg_8_ ( .D(n5384), .CK(clk), .QN(n4581) );
  DLH_X1 round_in_data_reg_8_ ( .G(n5471), .D(U49_Z_8), .Q(n3528) );
  DFF_X1 cipher_text_reg_8_ ( .D(n5385), .CK(clk), .Q(out_data[8]) );
  DFF_X1 temp_round_data_reg_9_ ( .D(n5382), .CK(clk), .QN(n4580) );
  DLH_X1 round_in_data_reg_9_ ( .G(n5471), .D(U49_Z_9), .Q(n3529) );
  DFF_X1 cipher_text_reg_9_ ( .D(n5383), .CK(clk), .Q(out_data[9]) );
  DFF_X1 temp_round_data_reg_10_ ( .D(n5380), .CK(clk), .QN(n4579) );
  DLH_X1 round_in_data_reg_10_ ( .G(U46_Z_1), .D(U49_Z_10), .Q(n3530) );
  DFF_X1 cipher_text_reg_10_ ( .D(n5381), .CK(clk), .Q(out_data[10]) );
  DFF_X1 temp_round_data_reg_11_ ( .D(n5378), .CK(clk), .QN(n4578) );
  DLH_X1 round_in_data_reg_11_ ( .G(U46_Z_1), .D(U49_Z_11), .Q(n3531) );
  DFF_X1 cipher_text_reg_11_ ( .D(n5379), .CK(clk), .Q(out_data[11]) );
  DFF_X1 temp_round_data_reg_12_ ( .D(n5376), .CK(clk), .QN(n4577) );
  DLH_X1 round_in_data_reg_12_ ( .G(n5471), .D(U49_Z_12), .Q(n3532) );
  DFF_X1 cipher_text_reg_12_ ( .D(n5377), .CK(clk), .Q(out_data[12]) );
  DFF_X1 temp_round_data_reg_13_ ( .D(n5374), .CK(clk), .QN(n4576) );
  DLH_X1 round_in_data_reg_13_ ( .G(n5464), .D(U49_Z_13), .Q(n3533) );
  DFF_X1 cipher_text_reg_13_ ( .D(n5375), .CK(clk), .Q(out_data[13]) );
  DFF_X1 temp_round_data_reg_14_ ( .D(n5372), .CK(clk), .QN(n4575) );
  DLH_X1 round_in_data_reg_14_ ( .G(n5465), .D(U49_Z_14), .Q(n3534) );
  DFF_X1 cipher_text_reg_14_ ( .D(n5373), .CK(clk), .Q(out_data[14]) );
  DFF_X1 temp_round_data_reg_15_ ( .D(n5370), .CK(clk), .QN(n4574) );
  DLH_X1 round_in_data_reg_15_ ( .G(n5470), .D(U49_Z_15), .Q(n3535) );
  DFF_X1 cipher_text_reg_15_ ( .D(n5371), .CK(clk), .Q(out_data[15]) );
  DFF_X1 temp_round_data_reg_16_ ( .D(n5368), .CK(clk), .QN(n4573) );
  DLH_X1 round_in_data_reg_16_ ( .G(U46_Z_1), .D(U49_Z_16), .Q(n3536) );
  DFF_X1 cipher_text_reg_16_ ( .D(n5369), .CK(clk), .Q(out_data[16]) );
  DFF_X1 temp_round_data_reg_17_ ( .D(n5366), .CK(clk), .QN(n4572) );
  DLH_X1 round_in_data_reg_17_ ( .G(n5468), .D(U49_Z_17), .Q(n3537) );
  DFF_X1 cipher_text_reg_17_ ( .D(n5367), .CK(clk), .Q(out_data[17]) );
  DFF_X1 temp_round_data_reg_18_ ( .D(n5364), .CK(clk), .QN(n4571) );
  DLH_X1 round_in_data_reg_18_ ( .G(n5470), .D(U49_Z_18), .Q(n3538) );
  DFF_X1 cipher_text_reg_18_ ( .D(n5365), .CK(clk), .Q(out_data[18]) );
  DFF_X1 temp_round_data_reg_19_ ( .D(n5362), .CK(clk), .QN(n4570) );
  DLH_X1 round_in_data_reg_19_ ( .G(n5469), .D(U49_Z_19), .Q(n3539) );
  DFF_X1 cipher_text_reg_19_ ( .D(n5363), .CK(clk), .Q(out_data[19]) );
  DFF_X1 temp_round_data_reg_20_ ( .D(n5360), .CK(clk), .QN(n4569) );
  DLH_X1 round_in_data_reg_20_ ( .G(n5467), .D(U49_Z_20), .Q(n3540) );
  DFF_X1 cipher_text_reg_20_ ( .D(n5361), .CK(clk), .Q(out_data[20]) );
  DFF_X1 temp_round_data_reg_21_ ( .D(n5358), .CK(clk), .QN(n4568) );
  DLH_X1 round_in_data_reg_21_ ( .G(n5471), .D(U49_Z_21), .Q(n3541) );
  DFF_X1 cipher_text_reg_21_ ( .D(n5359), .CK(clk), .Q(out_data[21]) );
  DFF_X1 temp_round_data_reg_22_ ( .D(n5356), .CK(clk), .QN(n4567) );
  DLH_X1 round_in_data_reg_22_ ( .G(n5465), .D(U49_Z_22), .Q(n3542) );
  DFF_X1 cipher_text_reg_22_ ( .D(n5357), .CK(clk), .Q(out_data[22]) );
  DFF_X1 temp_round_data_reg_23_ ( .D(n5354), .CK(clk), .QN(n4566) );
  DLH_X1 round_in_data_reg_23_ ( .G(n5464), .D(U49_Z_23), .Q(n3543) );
  DFF_X1 cipher_text_reg_23_ ( .D(n5355), .CK(clk), .Q(out_data[23]) );
  DFF_X1 temp_round_data_reg_24_ ( .D(n5352), .CK(clk), .QN(n4565) );
  DLH_X1 round_in_data_reg_24_ ( .G(n5469), .D(U49_Z_24), .Q(n3544) );
  DFF_X1 cipher_text_reg_24_ ( .D(n5353), .CK(clk), .Q(out_data[24]) );
  DFF_X1 temp_round_data_reg_25_ ( .D(n5350), .CK(clk), .QN(n4564) );
  DLH_X1 round_in_data_reg_25_ ( .G(n5466), .D(U49_Z_25), .Q(n3545) );
  DFF_X1 cipher_text_reg_25_ ( .D(n5351), .CK(clk), .Q(out_data[25]) );
  DFF_X1 temp_round_data_reg_26_ ( .D(n5348), .CK(clk), .QN(n4563) );
  DLH_X1 round_in_data_reg_26_ ( .G(n5465), .D(U49_Z_26), .Q(n3546) );
  DFF_X1 cipher_text_reg_26_ ( .D(n5349), .CK(clk), .Q(out_data[26]) );
  DFF_X1 temp_round_data_reg_27_ ( .D(n5346), .CK(clk), .QN(n4562) );
  DLH_X1 round_in_data_reg_27_ ( .G(n5470), .D(U49_Z_27), .Q(n3547) );
  DFF_X1 cipher_text_reg_27_ ( .D(n5347), .CK(clk), .Q(out_data[27]) );
  DFF_X1 temp_round_data_reg_28_ ( .D(n5344), .CK(clk), .QN(n4561) );
  DLH_X1 round_in_data_reg_28_ ( .G(n5464), .D(U49_Z_28), .Q(n3548) );
  DFF_X1 cipher_text_reg_28_ ( .D(n5345), .CK(clk), .Q(out_data[28]) );
  DFF_X1 temp_round_data_reg_29_ ( .D(n5342), .CK(clk), .QN(n4560) );
  DLH_X1 round_in_data_reg_29_ ( .G(n5471), .D(U49_Z_29), .Q(n3549) );
  DFF_X1 cipher_text_reg_29_ ( .D(n5343), .CK(clk), .Q(out_data[29]) );
  DFF_X1 temp_round_data_reg_30_ ( .D(n5340), .CK(clk), .QN(n4559) );
  DLH_X1 round_in_data_reg_30_ ( .G(n5470), .D(U49_Z_30), .Q(n3550) );
  DFF_X1 cipher_text_reg_30_ ( .D(n5341), .CK(clk), .Q(out_data[30]) );
  DFF_X1 temp_round_data_reg_31_ ( .D(n5338), .CK(clk), .QN(n4558) );
  DLH_X1 round_in_data_reg_31_ ( .G(n5468), .D(U49_Z_31), .Q(n3551) );
  DFF_X1 cipher_text_reg_31_ ( .D(n5339), .CK(clk), .Q(out_data[31]) );
  DFF_X1 temp_round_data_reg_32_ ( .D(n5336), .CK(clk), .QN(n4557) );
  DLH_X1 round_in_data_reg_32_ ( .G(n5469), .D(U49_Z_32), .Q(n3552) );
  DFF_X1 cipher_text_reg_32_ ( .D(n5337), .CK(clk), .Q(out_data[32]) );
  DFF_X1 temp_round_data_reg_33_ ( .D(n5334), .CK(clk), .QN(n4556) );
  DLH_X1 round_in_data_reg_33_ ( .G(n5470), .D(U49_Z_33), .Q(n3553) );
  DFF_X1 cipher_text_reg_33_ ( .D(n5335), .CK(clk), .Q(out_data[33]) );
  DFF_X1 temp_round_data_reg_34_ ( .D(n5332), .CK(clk), .QN(n4555) );
  DLH_X1 round_in_data_reg_34_ ( .G(n5465), .D(U49_Z_34), .Q(n3554) );
  DFF_X1 cipher_text_reg_34_ ( .D(n5333), .CK(clk), .Q(out_data[34]) );
  DFF_X1 temp_round_data_reg_35_ ( .D(n5330), .CK(clk), .QN(n4554) );
  DLH_X1 round_in_data_reg_35_ ( .G(n5469), .D(U49_Z_35), .Q(n3555) );
  DFF_X1 cipher_text_reg_35_ ( .D(n5331), .CK(clk), .Q(out_data[35]) );
  DFF_X1 temp_round_data_reg_36_ ( .D(n5328), .CK(clk), .QN(n4553) );
  DLH_X1 round_in_data_reg_36_ ( .G(n5467), .D(U49_Z_36), .Q(n3556) );
  DFF_X1 cipher_text_reg_36_ ( .D(n5329), .CK(clk), .Q(out_data[36]) );
  DFF_X1 temp_round_data_reg_37_ ( .D(n5326), .CK(clk), .QN(n4552) );
  DLH_X1 round_in_data_reg_37_ ( .G(n5466), .D(U49_Z_37), .Q(n3557) );
  DFF_X1 cipher_text_reg_37_ ( .D(n5327), .CK(clk), .Q(out_data[37]) );
  DFF_X1 temp_round_data_reg_38_ ( .D(n5324), .CK(clk), .QN(n4551) );
  DLH_X1 round_in_data_reg_38_ ( .G(n5468), .D(U49_Z_38), .Q(n3558) );
  DFF_X1 cipher_text_reg_38_ ( .D(n5325), .CK(clk), .Q(out_data[38]) );
  DFF_X1 temp_round_data_reg_39_ ( .D(n5322), .CK(clk), .QN(n4550) );
  DLH_X1 round_in_data_reg_39_ ( .G(n5467), .D(U49_Z_39), .Q(n3559) );
  DFF_X1 cipher_text_reg_39_ ( .D(n5323), .CK(clk), .Q(out_data[39]) );
  DFF_X1 temp_round_data_reg_40_ ( .D(n5320), .CK(clk), .QN(n4549) );
  DLH_X1 round_in_data_reg_40_ ( .G(n5471), .D(U49_Z_40), .Q(n3560) );
  DFF_X1 cipher_text_reg_40_ ( .D(n5321), .CK(clk), .Q(out_data[40]) );
  DFF_X1 temp_round_data_reg_41_ ( .D(n5318), .CK(clk), .QN(n4548) );
  DLH_X1 round_in_data_reg_41_ ( .G(n5468), .D(U49_Z_41), .Q(n3561) );
  DFF_X1 cipher_text_reg_41_ ( .D(n5319), .CK(clk), .Q(out_data[41]) );
  DFF_X1 temp_round_data_reg_42_ ( .D(n5316), .CK(clk), .QN(n4547) );
  DLH_X1 round_in_data_reg_42_ ( .G(n5465), .D(U49_Z_42), .Q(n3562) );
  DFF_X1 cipher_text_reg_42_ ( .D(n5317), .CK(clk), .Q(out_data[42]) );
  DFF_X1 temp_round_data_reg_43_ ( .D(n5314), .CK(clk), .QN(n4546) );
  DLH_X1 round_in_data_reg_43_ ( .G(n5470), .D(U49_Z_43), .Q(n3563) );
  DFF_X1 cipher_text_reg_43_ ( .D(n5315), .CK(clk), .Q(out_data[43]) );
  DFF_X1 temp_round_data_reg_44_ ( .D(n5312), .CK(clk), .QN(n4545) );
  DLH_X1 round_in_data_reg_44_ ( .G(n5464), .D(U49_Z_44), .Q(n3564) );
  DFF_X1 cipher_text_reg_44_ ( .D(n5313), .CK(clk), .Q(out_data[44]) );
  DFF_X1 temp_round_data_reg_45_ ( .D(n5310), .CK(clk), .QN(n4544) );
  DLH_X1 round_in_data_reg_45_ ( .G(n5464), .D(U49_Z_45), .Q(n3565) );
  DFF_X1 cipher_text_reg_45_ ( .D(n5311), .CK(clk), .Q(out_data[45]) );
  DFF_X1 temp_round_data_reg_46_ ( .D(n5308), .CK(clk), .QN(n4543) );
  DLH_X1 round_in_data_reg_46_ ( .G(n5466), .D(U49_Z_46), .Q(n3566) );
  DFF_X1 cipher_text_reg_46_ ( .D(n5309), .CK(clk), .Q(out_data[46]) );
  DFF_X1 temp_round_data_reg_47_ ( .D(n5306), .CK(clk), .QN(n4542) );
  DLH_X1 round_in_data_reg_47_ ( .G(n5466), .D(U49_Z_47), .Q(n3567) );
  DFF_X1 cipher_text_reg_47_ ( .D(n5307), .CK(clk), .Q(out_data[47]) );
  DFF_X1 temp_round_data_reg_48_ ( .D(n5304), .CK(clk), .QN(n4541) );
  DLH_X1 round_in_data_reg_48_ ( .G(n5464), .D(U49_Z_48), .Q(n3568) );
  DFF_X1 cipher_text_reg_48_ ( .D(n5305), .CK(clk), .Q(out_data[48]) );
  DFF_X1 temp_round_data_reg_49_ ( .D(n5302), .CK(clk), .QN(n4540) );
  DLH_X1 round_in_data_reg_49_ ( .G(n5469), .D(U49_Z_49), .Q(n3569) );
  DFF_X1 cipher_text_reg_49_ ( .D(n5303), .CK(clk), .Q(out_data[49]) );
  DFF_X1 temp_round_data_reg_50_ ( .D(n5300), .CK(clk), .QN(n4539) );
  DLH_X1 round_in_data_reg_50_ ( .G(n5469), .D(U49_Z_50), .Q(n3570) );
  DFF_X1 cipher_text_reg_50_ ( .D(n5301), .CK(clk), .Q(out_data[50]) );
  DFF_X1 temp_round_data_reg_51_ ( .D(n5298), .CK(clk), .QN(n4538) );
  DLH_X1 round_in_data_reg_51_ ( .G(n5465), .D(U49_Z_51), .Q(n3571) );
  DFF_X1 cipher_text_reg_51_ ( .D(n5299), .CK(clk), .Q(out_data[51]) );
  DFF_X1 temp_round_data_reg_52_ ( .D(n5296), .CK(clk), .QN(n4537) );
  DLH_X1 round_in_data_reg_52_ ( .G(n5471), .D(U49_Z_52), .Q(n3572) );
  DFF_X1 cipher_text_reg_52_ ( .D(n5297), .CK(clk), .Q(out_data[52]) );
  DFF_X1 temp_round_data_reg_53_ ( .D(n5294), .CK(clk), .QN(n4536) );
  DLH_X1 round_in_data_reg_53_ ( .G(n5465), .D(U49_Z_53), .Q(n3573) );
  DFF_X1 cipher_text_reg_53_ ( .D(n5295), .CK(clk), .Q(out_data[53]) );
  DFF_X1 temp_round_data_reg_54_ ( .D(n5292), .CK(clk), .QN(n4535) );
  DLH_X1 round_in_data_reg_54_ ( .G(n5470), .D(U49_Z_54), .Q(n3574) );
  DFF_X1 cipher_text_reg_54_ ( .D(n5293), .CK(clk), .Q(out_data[54]) );
  DFF_X1 temp_round_data_reg_55_ ( .D(n5290), .CK(clk), .QN(n4534) );
  DLH_X1 round_in_data_reg_55_ ( .G(n5470), .D(U49_Z_55), .Q(n3575) );
  DFF_X1 cipher_text_reg_55_ ( .D(n5291), .CK(clk), .Q(out_data[55]) );
  DFF_X1 temp_round_data_reg_56_ ( .D(n5288), .CK(clk), .QN(n4533) );
  DLH_X1 round_in_data_reg_56_ ( .G(n5471), .D(U49_Z_56), .Q(n3576) );
  DFF_X1 cipher_text_reg_56_ ( .D(n5289), .CK(clk), .Q(out_data[56]) );
  DFF_X1 temp_round_data_reg_57_ ( .D(n5286), .CK(clk), .QN(n4532) );
  DLH_X1 round_in_data_reg_57_ ( .G(n5467), .D(U49_Z_57), .Q(n3577) );
  DFF_X1 cipher_text_reg_57_ ( .D(n5287), .CK(clk), .Q(out_data[57]) );
  DFF_X1 temp_round_data_reg_58_ ( .D(n5284), .CK(clk), .QN(n4531) );
  DLH_X1 round_in_data_reg_58_ ( .G(n5468), .D(U49_Z_58), .Q(n3578) );
  DFF_X1 cipher_text_reg_58_ ( .D(n5285), .CK(clk), .Q(out_data[58]) );
  DFF_X1 temp_round_data_reg_59_ ( .D(n5282), .CK(clk), .QN(n4530) );
  DLH_X1 round_in_data_reg_59_ ( .G(n5464), .D(U49_Z_59), .Q(n3579) );
  DFF_X1 cipher_text_reg_59_ ( .D(n5283), .CK(clk), .Q(out_data[59]) );
  DFF_X1 temp_round_data_reg_60_ ( .D(n5280), .CK(clk), .QN(n4529) );
  DLH_X1 round_in_data_reg_60_ ( .G(n5466), .D(U49_Z_60), .Q(n3580) );
  DFF_X1 cipher_text_reg_60_ ( .D(n5281), .CK(clk), .Q(out_data[60]) );
  DFF_X1 temp_round_data_reg_61_ ( .D(n5278), .CK(clk), .QN(n4528) );
  DLH_X1 round_in_data_reg_61_ ( .G(n5471), .D(U49_Z_61), .Q(n3581) );
  DFF_X1 cipher_text_reg_61_ ( .D(n5279), .CK(clk), .Q(out_data[61]) );
  DFF_X1 temp_round_data_reg_62_ ( .D(n5276), .CK(clk), .QN(n4527) );
  DLH_X1 round_in_data_reg_62_ ( .G(U46_Z_1), .D(U49_Z_62), .Q(n3582) );
  DFF_X1 cipher_text_reg_62_ ( .D(n5277), .CK(clk), .Q(out_data[62]) );
  DFF_X1 temp_round_data_reg_63_ ( .D(n5274), .CK(clk), .QN(n4526) );
  DLH_X1 round_in_data_reg_63_ ( .G(n5471), .D(U49_Z_63), .Q(n3583) );
  DFF_X1 cipher_text_reg_63_ ( .D(n5275), .CK(clk), .Q(out_data[63]) );
  DFF_X1 temp_round_data_reg_64_ ( .D(n5272), .CK(clk), .QN(n4525) );
  DLH_X1 round_in_data_reg_64_ ( .G(n5471), .D(U49_Z_64), .Q(n3584) );
  DFF_X1 cipher_text_reg_64_ ( .D(n5273), .CK(clk), .Q(out_data[64]) );
  DFF_X1 temp_round_data_reg_65_ ( .D(n5270), .CK(clk), .QN(n4524) );
  DLH_X1 round_in_data_reg_65_ ( .G(n5465), .D(U49_Z_65), .Q(n3585) );
  DFF_X1 cipher_text_reg_65_ ( .D(n5271), .CK(clk), .Q(out_data[65]) );
  DFF_X1 temp_round_data_reg_66_ ( .D(n5268), .CK(clk), .QN(n4523) );
  DLH_X1 round_in_data_reg_66_ ( .G(U46_Z_1), .D(U49_Z_66), .Q(n3586) );
  DFF_X1 cipher_text_reg_66_ ( .D(n5269), .CK(clk), .Q(out_data[66]) );
  DFF_X1 temp_round_data_reg_67_ ( .D(n5266), .CK(clk), .QN(n4522) );
  DLH_X1 round_in_data_reg_67_ ( .G(n5471), .D(U49_Z_67), .Q(n3587) );
  DFF_X1 cipher_text_reg_67_ ( .D(n5267), .CK(clk), .Q(out_data[67]) );
  DFF_X1 temp_round_data_reg_68_ ( .D(n5264), .CK(clk), .QN(n4521) );
  DLH_X1 round_in_data_reg_68_ ( .G(n5471), .D(U49_Z_68), .Q(n3588) );
  DFF_X1 cipher_text_reg_68_ ( .D(n5265), .CK(clk), .Q(out_data[68]) );
  DFF_X1 temp_round_data_reg_69_ ( .D(n5262), .CK(clk), .QN(n4520) );
  DLH_X1 round_in_data_reg_69_ ( .G(n5469), .D(U49_Z_69), .Q(n3589) );
  DFF_X1 cipher_text_reg_69_ ( .D(n5263), .CK(clk), .Q(out_data[69]) );
  DFF_X1 temp_round_data_reg_70_ ( .D(n5260), .CK(clk), .QN(n4519) );
  DLH_X1 round_in_data_reg_70_ ( .G(n5471), .D(U49_Z_70), .Q(n3590) );
  DFF_X1 cipher_text_reg_70_ ( .D(n5261), .CK(clk), .Q(out_data[70]) );
  DFF_X1 temp_round_data_reg_71_ ( .D(n5258), .CK(clk), .QN(n4518) );
  DLH_X1 round_in_data_reg_71_ ( .G(n5467), .D(U49_Z_71), .Q(n3591) );
  DFF_X1 cipher_text_reg_71_ ( .D(n5259), .CK(clk), .Q(out_data[71]) );
  DFF_X1 temp_round_data_reg_72_ ( .D(n5256), .CK(clk), .QN(n4517) );
  DLH_X1 round_in_data_reg_72_ ( .G(n5464), .D(U49_Z_72), .Q(n3592) );
  DFF_X1 cipher_text_reg_72_ ( .D(n5257), .CK(clk), .Q(out_data[72]) );
  DFF_X1 temp_round_data_reg_73_ ( .D(n5254), .CK(clk), .QN(n4516) );
  DLH_X1 round_in_data_reg_73_ ( .G(n5468), .D(U49_Z_73), .Q(n3593) );
  DFF_X1 cipher_text_reg_73_ ( .D(n5255), .CK(clk), .Q(out_data[73]) );
  DFF_X1 temp_round_data_reg_74_ ( .D(n5252), .CK(clk), .QN(n4515) );
  DLH_X1 round_in_data_reg_74_ ( .G(n5466), .D(U49_Z_74), .Q(n3594) );
  DFF_X1 cipher_text_reg_74_ ( .D(n5253), .CK(clk), .Q(out_data[74]) );
  DFF_X1 temp_round_data_reg_75_ ( .D(n5250), .CK(clk), .QN(n4514) );
  DLH_X1 round_in_data_reg_75_ ( .G(n5470), .D(U49_Z_75), .Q(n3595) );
  DFF_X1 cipher_text_reg_75_ ( .D(n5251), .CK(clk), .Q(out_data[75]) );
  DFF_X1 temp_round_data_reg_76_ ( .D(n5248), .CK(clk), .QN(n4513) );
  DLH_X1 round_in_data_reg_76_ ( .G(n5469), .D(U49_Z_76), .Q(n3596) );
  DFF_X1 cipher_text_reg_76_ ( .D(n5249), .CK(clk), .Q(out_data[76]) );
  DFF_X1 temp_round_data_reg_77_ ( .D(n5246), .CK(clk), .QN(n4512) );
  DLH_X1 round_in_data_reg_77_ ( .G(n5466), .D(U49_Z_77), .Q(n3597) );
  DFF_X1 cipher_text_reg_77_ ( .D(n5247), .CK(clk), .Q(out_data[77]) );
  DFF_X1 temp_round_data_reg_78_ ( .D(n5244), .CK(clk), .QN(n4511) );
  DLH_X1 round_in_data_reg_78_ ( .G(n5470), .D(U49_Z_78), .Q(n3598) );
  DFF_X1 cipher_text_reg_78_ ( .D(n5245), .CK(clk), .Q(out_data[78]) );
  DFF_X1 temp_round_data_reg_79_ ( .D(n5242), .CK(clk), .QN(n4510) );
  DLH_X1 round_in_data_reg_79_ ( .G(n5469), .D(U49_Z_79), .Q(n3599) );
  DFF_X1 cipher_text_reg_79_ ( .D(n5243), .CK(clk), .Q(out_data[79]) );
  DFF_X1 temp_round_data_reg_80_ ( .D(n5240), .CK(clk), .QN(n4509) );
  DLH_X1 round_in_data_reg_80_ ( .G(n5467), .D(U49_Z_80), .Q(n3600) );
  DFF_X1 cipher_text_reg_80_ ( .D(n5241), .CK(clk), .Q(out_data[80]) );
  DFF_X1 temp_round_data_reg_81_ ( .D(n5238), .CK(clk), .QN(n4508) );
  DLH_X1 round_in_data_reg_81_ ( .G(n5471), .D(U49_Z_81), .Q(n3601) );
  DFF_X1 cipher_text_reg_81_ ( .D(n5239), .CK(clk), .Q(out_data[81]) );
  DFF_X1 temp_round_data_reg_82_ ( .D(n5236), .CK(clk), .QN(n4507) );
  DLH_X1 round_in_data_reg_82_ ( .G(n5465), .D(U49_Z_82), .Q(n3602) );
  DFF_X1 cipher_text_reg_82_ ( .D(n5237), .CK(clk), .Q(out_data[82]) );
  DFF_X1 temp_round_data_reg_83_ ( .D(n5234), .CK(clk), .QN(n4506) );
  DLH_X1 round_in_data_reg_83_ ( .G(U46_Z_1), .D(U49_Z_83), .Q(n3603) );
  DFF_X1 cipher_text_reg_83_ ( .D(n5235), .CK(clk), .Q(out_data[83]) );
  DFF_X1 temp_round_data_reg_84_ ( .D(n5232), .CK(clk), .QN(n4505) );
  DLH_X1 round_in_data_reg_84_ ( .G(n5468), .D(U49_Z_84), .Q(n3604) );
  DFF_X1 cipher_text_reg_84_ ( .D(n5233), .CK(clk), .Q(out_data[84]) );
  DFF_X1 temp_round_data_reg_85_ ( .D(n5230), .CK(clk), .QN(n4504) );
  DLH_X1 round_in_data_reg_85_ ( .G(n5468), .D(U49_Z_85), .Q(n3605) );
  DFF_X1 cipher_text_reg_85_ ( .D(n5231), .CK(clk), .Q(out_data[85]) );
  DFF_X1 temp_round_data_reg_86_ ( .D(n5228), .CK(clk), .QN(n4503) );
  DLH_X1 round_in_data_reg_86_ ( .G(n5471), .D(U49_Z_86), .Q(n3606) );
  DFF_X1 cipher_text_reg_86_ ( .D(n5229), .CK(clk), .Q(out_data[86]) );
  DFF_X1 temp_round_data_reg_87_ ( .D(n5226), .CK(clk), .QN(n4502) );
  DLH_X1 round_in_data_reg_87_ ( .G(n5468), .D(U49_Z_87), .Q(n3607) );
  DFF_X1 cipher_text_reg_87_ ( .D(n5227), .CK(clk), .Q(out_data[87]) );
  DFF_X1 temp_round_data_reg_88_ ( .D(n5224), .CK(clk), .QN(n4501) );
  DLH_X1 round_in_data_reg_88_ ( .G(n5469), .D(U49_Z_88), .Q(n3608) );
  DFF_X1 cipher_text_reg_88_ ( .D(n5225), .CK(clk), .Q(out_data[88]) );
  DFF_X1 temp_round_data_reg_89_ ( .D(n5222), .CK(clk), .QN(n4500) );
  DLH_X1 round_in_data_reg_89_ ( .G(n5465), .D(U49_Z_89), .Q(n3609) );
  DFF_X1 cipher_text_reg_89_ ( .D(n5223), .CK(clk), .Q(out_data[89]) );
  DFF_X1 temp_round_data_reg_90_ ( .D(n5220), .CK(clk), .QN(n4499) );
  DLH_X1 round_in_data_reg_90_ ( .G(n5471), .D(U49_Z_90), .Q(n3610) );
  DFF_X1 cipher_text_reg_90_ ( .D(n5221), .CK(clk), .Q(out_data[90]) );
  DFF_X1 temp_round_data_reg_91_ ( .D(n5218), .CK(clk), .QN(n4498) );
  DLH_X1 round_in_data_reg_91_ ( .G(n5471), .D(U49_Z_91), .Q(n3611) );
  DFF_X1 cipher_text_reg_91_ ( .D(n5219), .CK(clk), .Q(out_data[91]) );
  DFF_X1 temp_round_data_reg_92_ ( .D(n5216), .CK(clk), .QN(n4497) );
  DLH_X1 round_in_data_reg_92_ ( .G(n5466), .D(U49_Z_92), .Q(n3612) );
  DFF_X1 cipher_text_reg_92_ ( .D(n5217), .CK(clk), .Q(out_data[92]) );
  DFF_X1 temp_round_data_reg_93_ ( .D(n5214), .CK(clk), .QN(n4496) );
  DLH_X1 round_in_data_reg_93_ ( .G(n5465), .D(U49_Z_93), .Q(n3613) );
  DFF_X1 cipher_text_reg_93_ ( .D(n5215), .CK(clk), .Q(out_data[93]) );
  DFF_X1 temp_round_data_reg_94_ ( .D(n5212), .CK(clk), .QN(n4495) );
  DLH_X1 round_in_data_reg_94_ ( .G(n5470), .D(U49_Z_94), .Q(n3614) );
  DFF_X1 cipher_text_reg_94_ ( .D(n5213), .CK(clk), .Q(out_data[94]) );
  DFF_X1 temp_round_data_reg_95_ ( .D(n5210), .CK(clk), .QN(n4494) );
  DLH_X1 round_in_data_reg_95_ ( .G(n5467), .D(U49_Z_95), .Q(n3615) );
  DFF_X1 cipher_text_reg_95_ ( .D(n5211), .CK(clk), .Q(out_data[95]) );
  DFF_X1 temp_round_data_reg_96_ ( .D(n5208), .CK(clk), .QN(n4493) );
  DLH_X1 round_in_data_reg_96_ ( .G(n5464), .D(U49_Z_96), .Q(n3616) );
  DFF_X1 cipher_text_reg_96_ ( .D(n5209), .CK(clk), .Q(out_data[96]) );
  DFF_X1 temp_round_data_reg_97_ ( .D(n5206), .CK(clk), .QN(n4492) );
  DLH_X1 round_in_data_reg_97_ ( .G(n5467), .D(U49_Z_97), .Q(n3617) );
  DFF_X1 cipher_text_reg_97_ ( .D(n5207), .CK(clk), .Q(out_data[97]) );
  DFF_X1 temp_round_data_reg_98_ ( .D(n5204), .CK(clk), .QN(n4491) );
  DFF_X1 cipher_text_reg_98_ ( .D(n5205), .CK(clk), .Q(out_data[98]) );
  DFF_X1 temp_round_data_reg_99_ ( .D(n5202), .CK(clk), .QN(n4490) );
  DLH_X1 round_in_data_reg_99_ ( .G(n5464), .D(U49_Z_99), .Q(n3619) );
  DFF_X1 cipher_text_reg_99_ ( .D(n5203), .CK(clk), .Q(out_data[99]) );
  DFF_X1 temp_round_data_reg_100_ ( .D(n5200), .CK(clk), .QN(n4489) );
  DLH_X1 round_in_data_reg_100_ ( .G(n5468), .D(U49_Z_100), .Q(n3620) );
  DFF_X1 cipher_text_reg_100_ ( .D(n5201), .CK(clk), .Q(out_data[100]) );
  DFF_X1 temp_round_data_reg_101_ ( .D(n5198), .CK(clk), .QN(n4488) );
  DLH_X1 round_in_data_reg_101_ ( .G(n5469), .D(U49_Z_101), .Q(n3621) );
  DFF_X1 cipher_text_reg_101_ ( .D(n5199), .CK(clk), .Q(out_data[101]) );
  DFF_X1 temp_round_data_reg_102_ ( .D(n5196), .CK(clk), .QN(n4487) );
  DLH_X1 round_in_data_reg_102_ ( .G(n5469), .D(U49_Z_102), .Q(n3622) );
  DFF_X1 cipher_text_reg_102_ ( .D(n5197), .CK(clk), .Q(out_data[102]) );
  DFF_X1 temp_round_data_reg_103_ ( .D(n5194), .CK(clk), .QN(n4486) );
  DLH_X1 round_in_data_reg_103_ ( .G(n5466), .D(U49_Z_103), .Q(n3623) );
  DFF_X1 cipher_text_reg_103_ ( .D(n5195), .CK(clk), .Q(out_data[103]) );
  DFF_X1 temp_round_data_reg_104_ ( .D(n5192), .CK(clk), .QN(n4485) );
  DLH_X1 round_in_data_reg_104_ ( .G(n5466), .D(U49_Z_104), .Q(n3624) );
  DFF_X1 cipher_text_reg_104_ ( .D(n5193), .CK(clk), .Q(out_data[104]) );
  DFF_X1 temp_round_data_reg_105_ ( .D(n5190), .CK(clk), .QN(n4484) );
  DLH_X1 round_in_data_reg_105_ ( .G(n5465), .D(U49_Z_105), .Q(n3625) );
  DFF_X1 cipher_text_reg_105_ ( .D(n5191), .CK(clk), .Q(out_data[105]) );
  DFF_X1 temp_round_data_reg_106_ ( .D(n5188), .CK(clk), .QN(n4483) );
  DLH_X1 round_in_data_reg_106_ ( .G(n5467), .D(U49_Z_106), .Q(n3626) );
  DFF_X1 cipher_text_reg_106_ ( .D(n5189), .CK(clk), .Q(out_data[106]) );
  DFF_X1 temp_round_data_reg_107_ ( .D(n5186), .CK(clk), .QN(n4482) );
  DLH_X1 round_in_data_reg_107_ ( .G(n5465), .D(U49_Z_107), .Q(n3627) );
  DFF_X1 cipher_text_reg_107_ ( .D(n5187), .CK(clk), .Q(out_data[107]) );
  DFF_X1 temp_round_data_reg_108_ ( .D(n5184), .CK(clk), .QN(n4481) );
  DLH_X1 round_in_data_reg_108_ ( .G(n5469), .D(U49_Z_108), .Q(n3628) );
  DFF_X1 cipher_text_reg_108_ ( .D(n5185), .CK(clk), .Q(out_data[108]) );
  DFF_X1 temp_round_data_reg_109_ ( .D(n5182), .CK(clk), .QN(n4480) );
  DLH_X1 round_in_data_reg_109_ ( .G(n5466), .D(U49_Z_109), .Q(n3629) );
  DFF_X1 cipher_text_reg_109_ ( .D(n5183), .CK(clk), .Q(out_data[109]) );
  DFF_X1 temp_round_data_reg_110_ ( .D(n5180), .CK(clk), .QN(n4479) );
  DLH_X1 round_in_data_reg_110_ ( .G(n5470), .D(U49_Z_110), .Q(n3630) );
  DFF_X1 cipher_text_reg_110_ ( .D(n5181), .CK(clk), .Q(out_data[110]) );
  DFF_X1 temp_round_data_reg_111_ ( .D(n5178), .CK(clk), .QN(n4478) );
  DLH_X1 round_in_data_reg_111_ ( .G(n5467), .D(U49_Z_111), .Q(n3631) );
  DFF_X1 cipher_text_reg_111_ ( .D(n5179), .CK(clk), .Q(out_data[111]) );
  DFF_X1 temp_round_data_reg_112_ ( .D(n5176), .CK(clk), .QN(n4477) );
  DLH_X1 round_in_data_reg_112_ ( .G(n5466), .D(U49_Z_112), .Q(n3632) );
  DFF_X1 cipher_text_reg_112_ ( .D(n5177), .CK(clk), .Q(out_data[112]) );
  DFF_X1 temp_round_data_reg_113_ ( .D(n5174), .CK(clk), .QN(n4476) );
  DLH_X1 round_in_data_reg_113_ ( .G(U46_Z_1), .D(U49_Z_113), .Q(n3633) );
  DFF_X1 cipher_text_reg_113_ ( .D(n5175), .CK(clk), .Q(out_data[113]) );
  DFF_X1 temp_round_data_reg_114_ ( .D(n5172), .CK(clk), .QN(n4475) );
  DLH_X1 round_in_data_reg_114_ ( .G(n5468), .D(U49_Z_114), .Q(n3634) );
  DFF_X1 cipher_text_reg_114_ ( .D(n5173), .CK(clk), .Q(out_data[114]) );
  DFF_X1 temp_round_data_reg_115_ ( .D(n5170), .CK(clk), .QN(n4474) );
  DLH_X1 round_in_data_reg_115_ ( .G(n5464), .D(U49_Z_115), .Q(n3635) );
  DFF_X1 cipher_text_reg_115_ ( .D(n5171), .CK(clk), .Q(out_data[115]) );
  DFF_X1 temp_round_data_reg_116_ ( .D(n5168), .CK(clk), .QN(n4473) );
  DLH_X1 round_in_data_reg_116_ ( .G(n5464), .D(U49_Z_116), .Q(n3636) );
  DFF_X1 cipher_text_reg_116_ ( .D(n5169), .CK(clk), .Q(out_data[116]) );
  DFF_X1 temp_round_data_reg_117_ ( .D(n5166), .CK(clk), .QN(n4472) );
  DLH_X1 round_in_data_reg_117_ ( .G(U46_Z_1), .D(U49_Z_117), .Q(n3637) );
  DFF_X1 cipher_text_reg_117_ ( .D(n5167), .CK(clk), .Q(out_data[117]) );
  DFF_X1 temp_round_data_reg_118_ ( .D(n5164), .CK(clk), .QN(n4471) );
  DLH_X1 round_in_data_reg_118_ ( .G(n5471), .D(U49_Z_118), .Q(n3638) );
  DFF_X1 cipher_text_reg_118_ ( .D(n5165), .CK(clk), .Q(out_data[118]) );
  DFF_X1 temp_round_data_reg_119_ ( .D(n5162), .CK(clk), .QN(n4470) );
  DLH_X1 round_in_data_reg_119_ ( .G(n5471), .D(U49_Z_119), .Q(n3639) );
  DFF_X1 cipher_text_reg_119_ ( .D(n5163), .CK(clk), .Q(out_data[119]) );
  DFF_X1 temp_round_data_reg_120_ ( .D(n5160), .CK(clk), .QN(n4469) );
  DLH_X1 round_in_data_reg_120_ ( .G(n5471), .D(U49_Z_120), .Q(n3640) );
  DFF_X1 cipher_text_reg_120_ ( .D(n5161), .CK(clk), .Q(out_data[120]) );
  DFF_X1 temp_round_data_reg_121_ ( .D(n5158), .CK(clk), .QN(n4468) );
  DLH_X1 round_in_data_reg_121_ ( .G(n5464), .D(U49_Z_121), .Q(n3641) );
  DFF_X1 cipher_text_reg_121_ ( .D(n5159), .CK(clk), .Q(out_data[121]) );
  DFF_X1 temp_round_data_reg_122_ ( .D(n5156), .CK(clk), .QN(n4467) );
  DLH_X1 round_in_data_reg_122_ ( .G(n5464), .D(U49_Z_122), .Q(n3642) );
  DFF_X1 cipher_text_reg_122_ ( .D(n5157), .CK(clk), .Q(out_data[122]) );
  DFF_X1 temp_round_data_reg_123_ ( .D(n5154), .CK(clk), .QN(n4466) );
  DLH_X1 round_in_data_reg_123_ ( .G(U46_Z_1), .D(U49_Z_123), .Q(n3643) );
  DFF_X1 cipher_text_reg_123_ ( .D(n5155), .CK(clk), .Q(out_data[123]) );
  DFF_X1 temp_round_data_reg_124_ ( .D(n5152), .CK(clk), .QN(n4465) );
  DLH_X1 round_in_data_reg_124_ ( .G(n5467), .D(U49_Z_124), .Q(n3644) );
  DFF_X1 cipher_text_reg_124_ ( .D(n5153), .CK(clk), .Q(out_data[124]) );
  DFF_X1 temp_round_data_reg_125_ ( .D(n5150), .CK(clk), .QN(n4464) );
  DLH_X1 round_in_data_reg_125_ ( .G(U46_Z_1), .D(U49_Z_125), .Q(n3645) );
  DFF_X1 cipher_text_reg_125_ ( .D(n5151), .CK(clk), .Q(out_data[125]) );
  DFF_X1 temp_round_data_reg_126_ ( .D(n5148), .CK(clk), .QN(n4463) );
  DLH_X1 round_in_data_reg_126_ ( .G(n5470), .D(U49_Z_126), .Q(n3646) );
  DFF_X1 cipher_text_reg_126_ ( .D(n5149), .CK(clk), .Q(out_data[126]) );
  DFF_X1 temp_round_data_reg_127_ ( .D(n5146), .CK(clk), .QN(n4462) );
  DLH_X1 round_in_data_reg_127_ ( .G(U46_Z_1), .D(U49_Z_127), .Q(n3647) );
  DFF_X1 cipher_text_reg_127_ ( .D(n5147), .CK(clk), .Q(out_data[127]) );
  NAND3_X1 U1340 ( .A1(n5431), .A2(n4600), .A3(n4602), .ZN(n5405) );
  NAND4_X1 U1342 ( .A1(n4873), .A2(n4874), .A3(n4875), .A4(n4876), .ZN(n4870)
         );
  NAND3_X1 U1343 ( .A1(n4459), .A2(n5009), .A3(n4591), .ZN(U51_Z_1) );
  NAND3_X1 U1344 ( .A1(r424_A_1_), .A2(n5144), .A3(r424_A_2_), .ZN(n4866) );
  NAND3_X1 U1345 ( .A1(n4874), .A2(n4875), .A3(n4591), .ZN(U51_Z_2) );
  NAND3_X1 U1346 ( .A1(n5144), .A2(n4598), .A3(r424_A_2_), .ZN(n4873) );
  CLKBUF_X1 U1347 ( .A(U46_Z_1), .Z(n5464) );
  CLKBUF_X1 U1351 ( .A(n4601), .Z(n5453) );
  CLKBUF_X1 U1354 ( .A(n5431), .Z(n5442) );
  CLKBUF_X1 U1355 ( .A(n5442), .Z(n5440) );
  CLKBUF_X1 U1356 ( .A(n5442), .Z(n5439) );
  CLKBUF_X1 U1357 ( .A(n4602), .Z(n5445) );
  CLKBUF_X1 U1358 ( .A(n4602), .Z(n5444) );
  CLKBUF_X1 U1359 ( .A(n5444), .Z(n5452) );
  CLKBUF_X1 U1361 ( .A(n5443), .Z(n5446) );
  CLKBUF_X1 U1363 ( .A(n5445), .Z(n5450) );
  INV_X1 U1364 ( .A(n5431), .ZN(n5434) );
  INV_X1 U1365 ( .A(n5431), .ZN(n5435) );
  INV_X1 U1366 ( .A(n5442), .ZN(n5436) );
  INV_X1 U1367 ( .A(n5431), .ZN(n5437) );
  INV_X1 U1368 ( .A(n5442), .ZN(n5432) );
  INV_X1 U1369 ( .A(n5442), .ZN(n5433) );
  INV_X1 U1370 ( .A(n5463), .ZN(n5456) );
  INV_X1 U1371 ( .A(n5463), .ZN(n5455) );
  INV_X1 U1372 ( .A(n5430), .ZN(n5424) );
  INV_X1 U1373 ( .A(n5430), .ZN(n5422) );
  INV_X1 U1374 ( .A(n5427), .ZN(n5421) );
  INV_X1 U1375 ( .A(n5425), .ZN(n5423) );
  INV_X1 U1376 ( .A(n5419), .ZN(n5410) );
  INV_X1 U1377 ( .A(n5418), .ZN(n5409) );
  INV_X1 U1378 ( .A(n5419), .ZN(n5412) );
  INV_X1 U1379 ( .A(n5417), .ZN(n5413) );
  INV_X1 U1380 ( .A(n5419), .ZN(n5411) );
  BUF_X1 U1382 ( .A(n5442), .Z(n5438) );
  BUF_X1 U1383 ( .A(n5463), .Z(n5462) );
  BUF_X1 U1388 ( .A(n5416), .Z(n5414) );
  BUF_X1 U1389 ( .A(n5419), .Z(n5416) );
  BUF_X1 U1390 ( .A(n5430), .Z(n5426) );
  BUF_X1 U1391 ( .A(n5430), .Z(n5428) );
  BUF_X1 U1392 ( .A(n5430), .Z(n5427) );
  BUF_X1 U1393 ( .A(n5430), .Z(n5429) );
  INV_X1 U1394 ( .A(n5454), .ZN(n5463) );
  BUF_X1 U1395 ( .A(n5430), .Z(n5425) );
  INV_X1 U1396 ( .A(n5420), .ZN(n5430) );
  NOR3_X1 U1400 ( .A1(U51_Z_2), .A2(U51_Z_3), .A3(n5010), .ZN(n5143) );
  BUF_X1 U1401 ( .A(n4879), .Z(n5420) );
  NAND2_X1 U1402 ( .A1(n5405), .A2(n4600), .ZN(n4860) );
  INV_X1 U1403 ( .A(n5142), .ZN(n4595) );
  INV_X1 U1405 ( .A(n4865), .ZN(n4597) );
  NAND2_X1 U1406 ( .A1(n5144), .A2(n4595), .ZN(n4876) );
  NAND2_X1 U1407 ( .A1(n4865), .A2(n5144), .ZN(n4875) );
  INV_X1 U1408 ( .A(n4877), .ZN(n4592) );
  NAND2_X1 U1410 ( .A1(n5140), .A2(n4593), .ZN(n5012) );
  AND2_X1 U1411 ( .A1(n5008), .A2(n4872), .ZN(n5140) );
  NAND2_X1 U1412 ( .A1(n5007), .A2(n4872), .ZN(n4879) );
  AND2_X1 U1413 ( .A1(n5008), .A2(n4876), .ZN(n5007) );
  NAND2_X1 U1414 ( .A1(n4872), .A2(n4866), .ZN(U51_Z_3) );
  NAND2_X1 U1415 ( .A1(n4876), .A2(n5141), .ZN(n5010) );
  INV_X1 U1416 ( .A(n5408), .ZN(n4593) );
  INV_X1 U1417 ( .A(n5010), .ZN(n4459) );
  AND3_X1 U1418 ( .A1(n5141), .A2(n4590), .A3(n4866), .ZN(n5008) );
  INV_X1 U1419 ( .A(U51_Z_2), .ZN(n4590) );
  AND4_X1 U1420 ( .A1(n4875), .A2(n4873), .A3(n4866), .A4(n5009), .ZN(U51_Z_0)
         );
  NOR3_X1 U1421 ( .A1(rst), .A2(n3261), .A3(n2995), .ZN(n4730) );
  NOR3_X1 U1422 ( .A1(n4597), .A2(r424_A_0_), .A3(n4594), .ZN(n5408) );
  NOR2_X1 U1423 ( .A1(n4599), .A2(r424_A_3_), .ZN(n5144) );
  NOR2_X1 U1424 ( .A1(n4598), .A2(r424_A_2_), .ZN(n4865) );
  NOR2_X1 U1425 ( .A1(r424_A_0_), .A2(r424_A_3_), .ZN(n4877) );
  AOI21_X1 U1426 ( .B1(n4600), .B2(n4598), .A(n4862), .ZN(n4863) );
  OAI21_X1 U1427 ( .B1(rst), .B2(r424_A_0_), .A(n5405), .ZN(n4862) );
  INV_X1 U1428 ( .A(n4812), .ZN(n4119) );
  AOI22_X1 U1429 ( .A1(n5432), .A2(n[3048]), .B1(n5441), .B2(U99_DATA1_51), 
        .ZN(n4812) );
  INV_X1 U1430 ( .A(n4811), .ZN(n4120) );
  AOI22_X1 U1431 ( .A1(n5433), .A2(n[3047]), .B1(n5441), .B2(U99_DATA1_50), 
        .ZN(n4811) );
  INV_X1 U1432 ( .A(n4810), .ZN(n4121) );
  AOI22_X1 U1433 ( .A1(n5435), .A2(n[3046]), .B1(n5441), .B2(U99_DATA1_49), 
        .ZN(n4810) );
  INV_X1 U1434 ( .A(n4809), .ZN(n4122) );
  AOI22_X1 U1435 ( .A1(n5434), .A2(n[3045]), .B1(n5431), .B2(U99_DATA1_48), 
        .ZN(n4809) );
  INV_X1 U1436 ( .A(n4808), .ZN(n4123) );
  AOI22_X1 U1437 ( .A1(n5435), .A2(n[3044]), .B1(n5438), .B2(U99_DATA1_47), 
        .ZN(n4808) );
  INV_X1 U1438 ( .A(n4807), .ZN(n4124) );
  AOI22_X1 U1439 ( .A1(n5436), .A2(n[3043]), .B1(n5431), .B2(U99_DATA1_46), 
        .ZN(n4807) );
  INV_X1 U1440 ( .A(n4806), .ZN(n4125) );
  AOI22_X1 U1441 ( .A1(n5437), .A2(n[3042]), .B1(n5440), .B2(U99_DATA1_45), 
        .ZN(n4806) );
  INV_X1 U1442 ( .A(n4805), .ZN(n4126) );
  AOI22_X1 U1443 ( .A1(n5435), .A2(n[3041]), .B1(n5441), .B2(U99_DATA1_44), 
        .ZN(n4805) );
  OAI22_X1 U1444 ( .A1(n4860), .A2(n4866), .B1(n4863), .B2(n4594), .ZN(n5406)
         );
  OAI22_X1 U1445 ( .A1(n5457), .A2(n4326), .B1(n5458), .B2(n4465), .ZN(n5152)
         );
  OAI22_X1 U1446 ( .A1(n5457), .A2(n4325), .B1(n5463), .B2(n4466), .ZN(n5154)
         );
  OAI22_X1 U1447 ( .A1(n5457), .A2(n4324), .B1(n5461), .B2(n4467), .ZN(n5156)
         );
  OAI22_X1 U1448 ( .A1(n5457), .A2(n4323), .B1(n5459), .B2(n4468), .ZN(n5158)
         );
  OAI22_X1 U1449 ( .A1(n5457), .A2(n4322), .B1(n5462), .B2(n4469), .ZN(n5160)
         );
  OAI22_X1 U1450 ( .A1(n5454), .A2(n4321), .B1(n5458), .B2(n4470), .ZN(n5162)
         );
  OAI22_X1 U1451 ( .A1(n5454), .A2(n4320), .B1(n5459), .B2(n4471), .ZN(n5164)
         );
  OAI22_X1 U1452 ( .A1(n5454), .A2(n4319), .B1(n5458), .B2(n4472), .ZN(n5166)
         );
  OAI22_X1 U1453 ( .A1(n5454), .A2(n4318), .B1(n5458), .B2(n4473), .ZN(n5168)
         );
  OAI22_X1 U1454 ( .A1(n5456), .A2(n4317), .B1(n5461), .B2(n4474), .ZN(n5170)
         );
  OAI22_X1 U1455 ( .A1(n5455), .A2(n4316), .B1(n5461), .B2(n4475), .ZN(n5172)
         );
  OAI22_X1 U1456 ( .A1(n5453), .A2(n4315), .B1(n5460), .B2(n4476), .ZN(n5174)
         );
  OAI22_X1 U1457 ( .A1(n5454), .A2(n4314), .B1(n5461), .B2(n4477), .ZN(n5176)
         );
  OAI22_X1 U1458 ( .A1(n5455), .A2(n4313), .B1(n5461), .B2(n4478), .ZN(n5178)
         );
  OAI22_X1 U1459 ( .A1(n5453), .A2(n4312), .B1(n5459), .B2(n4479), .ZN(n5180)
         );
  OAI22_X1 U1460 ( .A1(n5456), .A2(n4311), .B1(n5463), .B2(n4480), .ZN(n5182)
         );
  OAI22_X1 U1461 ( .A1(n5454), .A2(n4310), .B1(n5459), .B2(n4481), .ZN(n5184)
         );
  OAI22_X1 U1462 ( .A1(n5456), .A2(n4309), .B1(n5462), .B2(n4482), .ZN(n5186)
         );
  OAI22_X1 U1463 ( .A1(n5456), .A2(n4308), .B1(n5461), .B2(n4483), .ZN(n5188)
         );
  OAI22_X1 U1464 ( .A1(n5455), .A2(n4307), .B1(n5463), .B2(n4484), .ZN(n5190)
         );
  OAI22_X1 U1465 ( .A1(n5457), .A2(n4306), .B1(n5460), .B2(n4485), .ZN(n5192)
         );
  OAI22_X1 U1466 ( .A1(n5453), .A2(n4305), .B1(n5459), .B2(n4486), .ZN(n5194)
         );
  OAI22_X1 U1467 ( .A1(n5453), .A2(n4304), .B1(n5458), .B2(n4487), .ZN(n5196)
         );
  OAI22_X1 U1468 ( .A1(n5453), .A2(n4303), .B1(n5462), .B2(n4488), .ZN(n5198)
         );
  OAI22_X1 U1469 ( .A1(n5453), .A2(n4302), .B1(n5462), .B2(n4489), .ZN(n5200)
         );
  OAI22_X1 U1470 ( .A1(n4601), .A2(n4301), .B1(n5461), .B2(n4490), .ZN(n5202)
         );
  OAI22_X1 U1471 ( .A1(n4601), .A2(n4300), .B1(n5462), .B2(n4491), .ZN(n5204)
         );
  OAI22_X1 U1472 ( .A1(n4601), .A2(n4299), .B1(n5460), .B2(n4492), .ZN(n5206)
         );
  OAI22_X1 U1473 ( .A1(n4601), .A2(n4298), .B1(n5460), .B2(n4493), .ZN(n5208)
         );
  OAI22_X1 U1474 ( .A1(n5454), .A2(n4297), .B1(n5462), .B2(n4494), .ZN(n5210)
         );
  OAI22_X1 U1475 ( .A1(n5454), .A2(n4296), .B1(n5458), .B2(n4495), .ZN(n5212)
         );
  OAI22_X1 U1476 ( .A1(n5454), .A2(n4295), .B1(n5460), .B2(n4496), .ZN(n5214)
         );
  OAI22_X1 U1477 ( .A1(n5454), .A2(n4294), .B1(n5461), .B2(n4497), .ZN(n5216)
         );
  OAI22_X1 U1478 ( .A1(n5454), .A2(n4293), .B1(n5459), .B2(n4498), .ZN(n5218)
         );
  OAI22_X1 U1479 ( .A1(n5454), .A2(n4292), .B1(n5460), .B2(n4499), .ZN(n5220)
         );
  OAI22_X1 U1480 ( .A1(n5454), .A2(n4291), .B1(n5459), .B2(n4500), .ZN(n5222)
         );
  OAI22_X1 U1481 ( .A1(n5454), .A2(n4290), .B1(n5461), .B2(n4501), .ZN(n5224)
         );
  OAI22_X1 U1482 ( .A1(n5454), .A2(n4289), .B1(n5460), .B2(n4502), .ZN(n5226)
         );
  OAI22_X1 U1483 ( .A1(n5454), .A2(n4288), .B1(n5461), .B2(n4503), .ZN(n5228)
         );
  OAI22_X1 U1484 ( .A1(n5454), .A2(n4287), .B1(n5458), .B2(n4504), .ZN(n5230)
         );
  OAI22_X1 U1485 ( .A1(n5454), .A2(n4286), .B1(n5462), .B2(n4505), .ZN(n5232)
         );
  OAI22_X1 U1486 ( .A1(n5454), .A2(n4285), .B1(n5458), .B2(n4506), .ZN(n5234)
         );
  OAI22_X1 U1487 ( .A1(n5456), .A2(n4284), .B1(n5459), .B2(n4507), .ZN(n5236)
         );
  OAI22_X1 U1488 ( .A1(n5455), .A2(n4283), .B1(n5463), .B2(n4508), .ZN(n5238)
         );
  OAI22_X1 U1489 ( .A1(n5455), .A2(n4282), .B1(n5458), .B2(n4509), .ZN(n5240)
         );
  OAI22_X1 U1490 ( .A1(n4601), .A2(n4281), .B1(n5458), .B2(n4510), .ZN(n5242)
         );
  OAI22_X1 U1491 ( .A1(n5454), .A2(n4280), .B1(n5458), .B2(n4511), .ZN(n5244)
         );
  OAI22_X1 U1492 ( .A1(n5455), .A2(n4279), .B1(n5459), .B2(n4512), .ZN(n5246)
         );
  OAI22_X1 U1493 ( .A1(n5456), .A2(n4278), .B1(n5459), .B2(n4513), .ZN(n5248)
         );
  OAI22_X1 U1494 ( .A1(n5455), .A2(n4277), .B1(n5458), .B2(n4514), .ZN(n5250)
         );
  OAI22_X1 U1495 ( .A1(n5456), .A2(n4276), .B1(n5459), .B2(n4515), .ZN(n5252)
         );
  OAI22_X1 U1496 ( .A1(n4601), .A2(n4275), .B1(n5462), .B2(n4516), .ZN(n5254)
         );
  OAI22_X1 U1497 ( .A1(n4601), .A2(n4274), .B1(n5460), .B2(n4517), .ZN(n5256)
         );
  OAI22_X1 U1498 ( .A1(n5457), .A2(n4273), .B1(n5460), .B2(n4518), .ZN(n5258)
         );
  OAI22_X1 U1499 ( .A1(n5457), .A2(n4272), .B1(n5460), .B2(n4519), .ZN(n5260)
         );
  OAI22_X1 U1500 ( .A1(n5457), .A2(n4271), .B1(n5459), .B2(n4520), .ZN(n5262)
         );
  OAI22_X1 U1501 ( .A1(n5457), .A2(n4270), .B1(n5460), .B2(n4521), .ZN(n5264)
         );
  OAI22_X1 U1502 ( .A1(n4601), .A2(n4269), .B1(n5459), .B2(n4522), .ZN(n5266)
         );
  OAI22_X1 U1503 ( .A1(n4601), .A2(n4268), .B1(n5462), .B2(n4523), .ZN(n5268)
         );
  OAI22_X1 U1504 ( .A1(n5457), .A2(n4267), .B1(n5458), .B2(n4524), .ZN(n5270)
         );
  OAI22_X1 U1505 ( .A1(n5453), .A2(n4266), .B1(n5461), .B2(n4525), .ZN(n5272)
         );
  OAI22_X1 U1506 ( .A1(n5453), .A2(n4265), .B1(n5458), .B2(n4526), .ZN(n5274)
         );
  OAI22_X1 U1507 ( .A1(n5454), .A2(n4264), .B1(n5458), .B2(n4527), .ZN(n5276)
         );
  OAI22_X1 U1508 ( .A1(n4601), .A2(n4263), .B1(n5459), .B2(n4528), .ZN(n5278)
         );
  OAI22_X1 U1509 ( .A1(n4601), .A2(n4262), .B1(n5459), .B2(n4529), .ZN(n5280)
         );
  OAI22_X1 U1510 ( .A1(n5454), .A2(n4261), .B1(n5461), .B2(n4530), .ZN(n5282)
         );
  OAI22_X1 U1511 ( .A1(n4601), .A2(n4260), .B1(n5458), .B2(n4531), .ZN(n5284)
         );
  OAI22_X1 U1512 ( .A1(n4601), .A2(n4259), .B1(n5458), .B2(n4532), .ZN(n5286)
         );
  OAI22_X1 U1513 ( .A1(n5457), .A2(n4258), .B1(n5458), .B2(n4533), .ZN(n5288)
         );
  OAI22_X1 U1514 ( .A1(n5457), .A2(n4257), .B1(n5461), .B2(n4534), .ZN(n5290)
         );
  OAI22_X1 U1515 ( .A1(n5453), .A2(n4256), .B1(n5462), .B2(n4535), .ZN(n5292)
         );
  OAI22_X1 U1516 ( .A1(n5457), .A2(n4255), .B1(n5463), .B2(n4536), .ZN(n5294)
         );
  OAI22_X1 U1517 ( .A1(n4601), .A2(n4254), .B1(n5460), .B2(n4537), .ZN(n5296)
         );
  OAI22_X1 U1518 ( .A1(n5457), .A2(n4253), .B1(n5461), .B2(n4538), .ZN(n5298)
         );
  OAI22_X1 U1519 ( .A1(n4601), .A2(n4252), .B1(n5461), .B2(n4539), .ZN(n5300)
         );
  OAI22_X1 U1520 ( .A1(n4601), .A2(n4251), .B1(n5460), .B2(n4540), .ZN(n5302)
         );
  OAI22_X1 U1521 ( .A1(n4601), .A2(n4250), .B1(n5460), .B2(n4541), .ZN(n5304)
         );
  OAI22_X1 U1522 ( .A1(n4601), .A2(n4249), .B1(n5460), .B2(n4542), .ZN(n5306)
         );
  OAI22_X1 U1523 ( .A1(n4601), .A2(n4248), .B1(n5462), .B2(n4543), .ZN(n5308)
         );
  OAI22_X1 U1524 ( .A1(n5457), .A2(n4247), .B1(n5462), .B2(n4544), .ZN(n5310)
         );
  OAI22_X1 U1525 ( .A1(n5454), .A2(n4246), .B1(n5459), .B2(n4545), .ZN(n5312)
         );
  OAI22_X1 U1526 ( .A1(n4601), .A2(n4245), .B1(n5460), .B2(n4546), .ZN(n5314)
         );
  OAI22_X1 U1527 ( .A1(n5454), .A2(n4244), .B1(n5461), .B2(n4547), .ZN(n5316)
         );
  OAI22_X1 U1528 ( .A1(n5453), .A2(n4243), .B1(n5458), .B2(n4548), .ZN(n5318)
         );
  OAI22_X1 U1529 ( .A1(n4601), .A2(n4242), .B1(n5458), .B2(n4549), .ZN(n5320)
         );
  OAI22_X1 U1530 ( .A1(n5457), .A2(n4241), .B1(n5462), .B2(n4550), .ZN(n5322)
         );
  OAI22_X1 U1531 ( .A1(n5453), .A2(n4240), .B1(n5462), .B2(n4551), .ZN(n5324)
         );
  OAI22_X1 U1532 ( .A1(n4601), .A2(n4239), .B1(n5460), .B2(n4552), .ZN(n5326)
         );
  OAI22_X1 U1533 ( .A1(n4601), .A2(n4238), .B1(n5462), .B2(n4553), .ZN(n5328)
         );
  OAI22_X1 U1534 ( .A1(n5456), .A2(n4237), .B1(n5460), .B2(n4554), .ZN(n5330)
         );
  OAI22_X1 U1535 ( .A1(n5456), .A2(n4236), .B1(n5458), .B2(n4555), .ZN(n5332)
         );
  OAI22_X1 U1536 ( .A1(n5456), .A2(n4235), .B1(n5460), .B2(n4556), .ZN(n5334)
         );
  OAI22_X1 U1537 ( .A1(n5456), .A2(n4234), .B1(n5462), .B2(n4557), .ZN(n5336)
         );
  OAI22_X1 U1538 ( .A1(n5456), .A2(n4233), .B1(n5459), .B2(n4558), .ZN(n5338)
         );
  OAI22_X1 U1539 ( .A1(n5456), .A2(n4232), .B1(n5461), .B2(n4559), .ZN(n5340)
         );
  OAI22_X1 U1540 ( .A1(n5456), .A2(n4231), .B1(n5461), .B2(n4560), .ZN(n5342)
         );
  OAI22_X1 U1541 ( .A1(n5456), .A2(n4230), .B1(n5461), .B2(n4561), .ZN(n5344)
         );
  OAI22_X1 U1542 ( .A1(n5456), .A2(n4229), .B1(n5462), .B2(n4562), .ZN(n5346)
         );
  OAI22_X1 U1543 ( .A1(n5456), .A2(n4228), .B1(n5461), .B2(n4563), .ZN(n5348)
         );
  OAI22_X1 U1544 ( .A1(n5456), .A2(n4227), .B1(n5461), .B2(n4564), .ZN(n5350)
         );
  OAI22_X1 U1545 ( .A1(n5456), .A2(n4226), .B1(n5459), .B2(n4565), .ZN(n5352)
         );
  OAI22_X1 U1546 ( .A1(n5455), .A2(n4225), .B1(n5459), .B2(n4566), .ZN(n5354)
         );
  OAI22_X1 U1547 ( .A1(n5455), .A2(n4224), .B1(n5458), .B2(n4567), .ZN(n5356)
         );
  OAI22_X1 U1548 ( .A1(n5455), .A2(n4223), .B1(n5459), .B2(n4568), .ZN(n5358)
         );
  OAI22_X1 U1549 ( .A1(n5455), .A2(n4222), .B1(n5459), .B2(n4569), .ZN(n5360)
         );
  OAI22_X1 U1550 ( .A1(n5455), .A2(n4221), .B1(n5460), .B2(n4570), .ZN(n5362)
         );
  OAI22_X1 U1551 ( .A1(n5455), .A2(n4220), .B1(n5458), .B2(n4571), .ZN(n5364)
         );
  OAI22_X1 U1552 ( .A1(n5455), .A2(n4219), .B1(n5458), .B2(n4572), .ZN(n5366)
         );
  OAI22_X1 U1553 ( .A1(n5455), .A2(n4218), .B1(n5462), .B2(n4573), .ZN(n5368)
         );
  OAI22_X1 U1554 ( .A1(n5455), .A2(n4217), .B1(n5460), .B2(n4574), .ZN(n5370)
         );
  OAI22_X1 U1555 ( .A1(n5455), .A2(n4216), .B1(n5460), .B2(n4575), .ZN(n5372)
         );
  OAI22_X1 U1556 ( .A1(n5455), .A2(n4215), .B1(n5461), .B2(n4576), .ZN(n5374)
         );
  OAI22_X1 U1557 ( .A1(n5455), .A2(n4214), .B1(n5459), .B2(n4577), .ZN(n5376)
         );
  OAI22_X1 U1558 ( .A1(n5453), .A2(n4213), .B1(n5459), .B2(n4578), .ZN(n5378)
         );
  OAI22_X1 U1559 ( .A1(n5453), .A2(n4212), .B1(n5460), .B2(n4579), .ZN(n5380)
         );
  OAI22_X1 U1560 ( .A1(n5453), .A2(n4211), .B1(n5461), .B2(n4580), .ZN(n5382)
         );
  OAI22_X1 U1561 ( .A1(n5453), .A2(n4210), .B1(n5460), .B2(n4581), .ZN(n5384)
         );
  OAI22_X1 U1562 ( .A1(n5453), .A2(n4209), .B1(n5459), .B2(n4582), .ZN(n5386)
         );
  OAI22_X1 U1563 ( .A1(n5453), .A2(n4208), .B1(n5458), .B2(n4583), .ZN(n5388)
         );
  OAI22_X1 U1564 ( .A1(n5453), .A2(n4207), .B1(n5461), .B2(n4584), .ZN(n5390)
         );
  OAI22_X1 U1565 ( .A1(n5453), .A2(n4206), .B1(n5459), .B2(n4585), .ZN(n5392)
         );
  OAI22_X1 U1566 ( .A1(n5453), .A2(n4205), .B1(n5460), .B2(n4586), .ZN(n5394)
         );
  OAI22_X1 U1567 ( .A1(n5453), .A2(n4204), .B1(n5462), .B2(n4587), .ZN(n5396)
         );
  OAI22_X1 U1568 ( .A1(n5453), .A2(n4203), .B1(n5461), .B2(n4588), .ZN(n5398)
         );
  OAI22_X1 U1569 ( .A1(n5453), .A2(n4202), .B1(n5461), .B2(n4589), .ZN(n5400)
         );
  OAI22_X1 U1570 ( .A1(n4863), .A2(n4596), .B1(n4860), .B2(n4864), .ZN(n5404)
         );
  NAND2_X1 U1571 ( .A1(n4865), .A2(r424_A_0_), .ZN(n4864) );
  OAI22_X1 U1572 ( .A1(n4070), .A2(n4598), .B1(n4860), .B2(n4861), .ZN(n5403)
         );
  NAND2_X1 U1573 ( .A1(r424_A_0_), .A2(n4598), .ZN(n4861) );
  INV_X1 U1574 ( .A(n4862), .ZN(n4070) );
  OAI22_X1 U1575 ( .A1(n5457), .A2(n4329), .B1(n5458), .B2(n4462), .ZN(n5146)
         );
  OAI22_X1 U1576 ( .A1(n5457), .A2(n4328), .B1(n5460), .B2(n4463), .ZN(n5148)
         );
  OAI22_X1 U1577 ( .A1(n5457), .A2(n4327), .B1(n5459), .B2(n4464), .ZN(n5150)
         );
  OAI22_X1 U1578 ( .A1(n4599), .A2(n5405), .B1(r424_A_0_), .B2(n4860), .ZN(
        n5407) );
  NAND2_X1 U1579 ( .A1(r424_A_3_), .A2(n4595), .ZN(n4872) );
  AND3_X1 U1581 ( .A1(n2996), .A2(n4595), .A3(n4877), .ZN(n4868) );
  NAND2_X1 U1582 ( .A1(n4596), .A2(n4598), .ZN(n5142) );
  NAND2_X1 U1583 ( .A1(r424_A_2_), .A2(n4877), .ZN(n4874) );
  INV_X1 U1584 ( .A(n4869), .ZN(n4201) );
  OAI211_X1 U1585 ( .C1(n4870), .C2(n4871), .A(n2996), .B(n3262), .ZN(n4869)
         );
  OAI211_X1 U1586 ( .C1(n4597), .C2(n4592), .A(n4872), .B(n4866), .ZN(n4871)
         );
  INV_X1 U1587 ( .A(n4760), .ZN(n4171) );
  AOI22_X1 U1588 ( .A1(n5436), .A2(n[3123]), .B1(n5440), .B2(U99_DATA1_126), 
        .ZN(n4760) );
  INV_X1 U1589 ( .A(n4759), .ZN(n4172) );
  AOI22_X1 U1590 ( .A1(n5437), .A2(n[3122]), .B1(n5441), .B2(U99_DATA1_125), 
        .ZN(n4759) );
  INV_X1 U1591 ( .A(n4758), .ZN(n4173) );
  AOI22_X1 U1592 ( .A1(n5432), .A2(n[3121]), .B1(n5439), .B2(U99_DATA1_124), 
        .ZN(n4758) );
  INV_X1 U1593 ( .A(n4757), .ZN(n4174) );
  AOI22_X1 U1594 ( .A1(n5433), .A2(n[3120]), .B1(n5441), .B2(U99_DATA1_123), 
        .ZN(n4757) );
  INV_X1 U1595 ( .A(n4756), .ZN(n4175) );
  AOI22_X1 U1596 ( .A1(n5434), .A2(n[3119]), .B1(n5441), .B2(U99_DATA1_122), 
        .ZN(n4756) );
  INV_X1 U1597 ( .A(n4755), .ZN(n4176) );
  AOI22_X1 U1598 ( .A1(n5435), .A2(n[3118]), .B1(n5441), .B2(U99_DATA1_121), 
        .ZN(n4755) );
  INV_X1 U1599 ( .A(n4754), .ZN(n4177) );
  AOI22_X1 U1600 ( .A1(n5436), .A2(n[3117]), .B1(n5438), .B2(U99_DATA1_120), 
        .ZN(n4754) );
  INV_X1 U1601 ( .A(n4753), .ZN(n4178) );
  AOI22_X1 U1602 ( .A1(n5437), .A2(n[3116]), .B1(n5440), .B2(U99_DATA1_119), 
        .ZN(n4753) );
  INV_X1 U1603 ( .A(n4752), .ZN(n4179) );
  AOI22_X1 U1604 ( .A1(n5434), .A2(n[3115]), .B1(n5441), .B2(U99_DATA1_118), 
        .ZN(n4752) );
  INV_X1 U1605 ( .A(n4751), .ZN(n4180) );
  AOI22_X1 U1606 ( .A1(n5434), .A2(n[3114]), .B1(n5439), .B2(U99_DATA1_117), 
        .ZN(n4751) );
  INV_X1 U1607 ( .A(n4750), .ZN(n4181) );
  AOI22_X1 U1608 ( .A1(n5434), .A2(n[3113]), .B1(n5441), .B2(U99_DATA1_116), 
        .ZN(n4750) );
  INV_X1 U1609 ( .A(n4749), .ZN(n4182) );
  AOI22_X1 U1610 ( .A1(n5434), .A2(n[3112]), .B1(n5431), .B2(U99_DATA1_115), 
        .ZN(n4749) );
  INV_X1 U1611 ( .A(n4748), .ZN(n4183) );
  AOI22_X1 U1612 ( .A1(n5434), .A2(n[3111]), .B1(n5431), .B2(U99_DATA1_114), 
        .ZN(n4748) );
  INV_X1 U1613 ( .A(n4747), .ZN(n4184) );
  AOI22_X1 U1614 ( .A1(n5434), .A2(n[3110]), .B1(n5441), .B2(U99_DATA1_113), 
        .ZN(n4747) );
  INV_X1 U1615 ( .A(n4746), .ZN(n4185) );
  AOI22_X1 U1616 ( .A1(n5434), .A2(n[3109]), .B1(n5440), .B2(U99_DATA1_112), 
        .ZN(n4746) );
  INV_X1 U1617 ( .A(n4745), .ZN(n4186) );
  AOI22_X1 U1618 ( .A1(n5434), .A2(n[3108]), .B1(n5438), .B2(U99_DATA1_111), 
        .ZN(n4745) );
  INV_X1 U1619 ( .A(n4744), .ZN(n4187) );
  AOI22_X1 U1620 ( .A1(n5434), .A2(n[3107]), .B1(n5431), .B2(U99_DATA1_110), 
        .ZN(n4744) );
  INV_X1 U1621 ( .A(n4743), .ZN(n4188) );
  AOI22_X1 U1622 ( .A1(n5434), .A2(n[3106]), .B1(n4733), .B2(U99_DATA1_109), 
        .ZN(n4743) );
  INV_X1 U1623 ( .A(n4742), .ZN(n4189) );
  AOI22_X1 U1624 ( .A1(n5434), .A2(n[3105]), .B1(n4733), .B2(U99_DATA1_108), 
        .ZN(n4742) );
  INV_X1 U1625 ( .A(n4741), .ZN(n4190) );
  AOI22_X1 U1626 ( .A1(n5434), .A2(n[3104]), .B1(n5439), .B2(U99_DATA1_107), 
        .ZN(n4741) );
  INV_X1 U1627 ( .A(n4740), .ZN(n4191) );
  AOI22_X1 U1628 ( .A1(n5435), .A2(n[3103]), .B1(n5438), .B2(U99_DATA1_106), 
        .ZN(n4740) );
  INV_X1 U1629 ( .A(n4739), .ZN(n4192) );
  AOI22_X1 U1630 ( .A1(n5435), .A2(n[3102]), .B1(n5431), .B2(U99_DATA1_105), 
        .ZN(n4739) );
  INV_X1 U1631 ( .A(n4738), .ZN(n4193) );
  AOI22_X1 U1632 ( .A1(n5435), .A2(n[3101]), .B1(n5440), .B2(U99_DATA1_104), 
        .ZN(n4738) );
  INV_X1 U1633 ( .A(n4737), .ZN(n4194) );
  AOI22_X1 U1634 ( .A1(n5435), .A2(n[3100]), .B1(n4733), .B2(U99_DATA1_103), 
        .ZN(n4737) );
  INV_X1 U1635 ( .A(n4736), .ZN(n4195) );
  AOI22_X1 U1636 ( .A1(n5435), .A2(n[3099]), .B1(n4733), .B2(U99_DATA1_102), 
        .ZN(n4736) );
  INV_X1 U1637 ( .A(n4735), .ZN(n4196) );
  AOI22_X1 U1638 ( .A1(n5435), .A2(n[3098]), .B1(n5441), .B2(U99_DATA1_101), 
        .ZN(n4735) );
  INV_X1 U1639 ( .A(n4734), .ZN(n4197) );
  AOI22_X1 U1640 ( .A1(n5435), .A2(n[3097]), .B1(n5441), .B2(U99_DATA1_100), 
        .ZN(n4734) );
  INV_X1 U1641 ( .A(n4732), .ZN(n4198) );
  AOI22_X1 U1642 ( .A1(n5435), .A2(n[3096]), .B1(n5439), .B2(U99_DATA1_99), 
        .ZN(n4732) );
  INV_X1 U1643 ( .A(n4859), .ZN(n4072) );
  AOI22_X1 U1644 ( .A1(n5437), .A2(n[3095]), .B1(n5438), .B2(U99_DATA1_98), 
        .ZN(n4859) );
  INV_X1 U1645 ( .A(n4858), .ZN(n4073) );
  AOI22_X1 U1646 ( .A1(n5434), .A2(n[3094]), .B1(n5441), .B2(U99_DATA1_97), 
        .ZN(n4858) );
  INV_X1 U1647 ( .A(n4857), .ZN(n4074) );
  AOI22_X1 U1648 ( .A1(n5432), .A2(n[3093]), .B1(n5431), .B2(U99_DATA1_96), 
        .ZN(n4857) );
  INV_X1 U1649 ( .A(n4856), .ZN(n4075) );
  AOI22_X1 U1650 ( .A1(n5433), .A2(n[3092]), .B1(n5439), .B2(U99_DATA1_95), 
        .ZN(n4856) );
  INV_X1 U1651 ( .A(n4855), .ZN(n4076) );
  AOI22_X1 U1652 ( .A1(n5434), .A2(n[3091]), .B1(n4733), .B2(U99_DATA1_94), 
        .ZN(n4855) );
  INV_X1 U1653 ( .A(n4854), .ZN(n4077) );
  AOI22_X1 U1654 ( .A1(n5434), .A2(n[3090]), .B1(n4733), .B2(U99_DATA1_93), 
        .ZN(n4854) );
  INV_X1 U1655 ( .A(n4853), .ZN(n4078) );
  AOI22_X1 U1656 ( .A1(n5435), .A2(n[3089]), .B1(n5431), .B2(U99_DATA1_92), 
        .ZN(n4853) );
  INV_X1 U1657 ( .A(n4852), .ZN(n4079) );
  AOI22_X1 U1658 ( .A1(n5435), .A2(n[3088]), .B1(n4733), .B2(U99_DATA1_91), 
        .ZN(n4852) );
  INV_X1 U1659 ( .A(n4851), .ZN(n4080) );
  AOI22_X1 U1660 ( .A1(n5435), .A2(n[3087]), .B1(n5431), .B2(U99_DATA1_90), 
        .ZN(n4851) );
  INV_X1 U1661 ( .A(n4850), .ZN(n4081) );
  AOI22_X1 U1662 ( .A1(n5435), .A2(n[3086]), .B1(n5441), .B2(U99_DATA1_89), 
        .ZN(n4850) );
  INV_X1 U1663 ( .A(n4849), .ZN(n4082) );
  AOI22_X1 U1664 ( .A1(n5435), .A2(n[3085]), .B1(n5431), .B2(U99_DATA1_88), 
        .ZN(n4849) );
  INV_X1 U1665 ( .A(n4848), .ZN(n4083) );
  AOI22_X1 U1666 ( .A1(n5436), .A2(n[3084]), .B1(n5431), .B2(U99_DATA1_87), 
        .ZN(n4848) );
  INV_X1 U1667 ( .A(n4847), .ZN(n4084) );
  AOI22_X1 U1668 ( .A1(n5436), .A2(n[3083]), .B1(n5441), .B2(U99_DATA1_86), 
        .ZN(n4847) );
  INV_X1 U1669 ( .A(n4846), .ZN(n4085) );
  AOI22_X1 U1670 ( .A1(n5436), .A2(n[3082]), .B1(n5441), .B2(U99_DATA1_85), 
        .ZN(n4846) );
  INV_X1 U1671 ( .A(n4845), .ZN(n4086) );
  AOI22_X1 U1672 ( .A1(n5436), .A2(n[3081]), .B1(n5441), .B2(U99_DATA1_84), 
        .ZN(n4845) );
  INV_X1 U1673 ( .A(n4844), .ZN(n4087) );
  AOI22_X1 U1674 ( .A1(n5436), .A2(n[3080]), .B1(n5439), .B2(U99_DATA1_83), 
        .ZN(n4844) );
  INV_X1 U1675 ( .A(n4843), .ZN(n4088) );
  AOI22_X1 U1676 ( .A1(n5436), .A2(n[3079]), .B1(n5439), .B2(U99_DATA1_82), 
        .ZN(n4843) );
  INV_X1 U1677 ( .A(n4842), .ZN(n4089) );
  AOI22_X1 U1678 ( .A1(n5436), .A2(n[3078]), .B1(n5438), .B2(U99_DATA1_81), 
        .ZN(n4842) );
  INV_X1 U1679 ( .A(n4841), .ZN(n4090) );
  AOI22_X1 U1680 ( .A1(n5436), .A2(n[3077]), .B1(n5441), .B2(U99_DATA1_80), 
        .ZN(n4841) );
  INV_X1 U1681 ( .A(n4840), .ZN(n4091) );
  AOI22_X1 U1682 ( .A1(n5436), .A2(n[3076]), .B1(n5438), .B2(U99_DATA1_79), 
        .ZN(n4840) );
  INV_X1 U1683 ( .A(n4839), .ZN(n4092) );
  AOI22_X1 U1684 ( .A1(n5437), .A2(n[3075]), .B1(n5441), .B2(U99_DATA1_78), 
        .ZN(n4839) );
  INV_X1 U1685 ( .A(n4838), .ZN(n4093) );
  AOI22_X1 U1686 ( .A1(n5434), .A2(n[3074]), .B1(n5440), .B2(U99_DATA1_77), 
        .ZN(n4838) );
  INV_X1 U1687 ( .A(n4837), .ZN(n4094) );
  AOI22_X1 U1688 ( .A1(n5435), .A2(n[3073]), .B1(n5441), .B2(U99_DATA1_76), 
        .ZN(n4837) );
  INV_X1 U1689 ( .A(n4836), .ZN(n4095) );
  AOI22_X1 U1690 ( .A1(n5437), .A2(n[3072]), .B1(n5441), .B2(U99_DATA1_75), 
        .ZN(n4836) );
  INV_X1 U1691 ( .A(n4835), .ZN(n4096) );
  AOI22_X1 U1692 ( .A1(n5437), .A2(n[3071]), .B1(n5441), .B2(U99_DATA1_74), 
        .ZN(n4835) );
  INV_X1 U1693 ( .A(n4834), .ZN(n4097) );
  AOI22_X1 U1694 ( .A1(n5437), .A2(n[3070]), .B1(n5441), .B2(U99_DATA1_73), 
        .ZN(n4834) );
  INV_X1 U1695 ( .A(n4833), .ZN(n4098) );
  AOI22_X1 U1696 ( .A1(n5437), .A2(n[3069]), .B1(n5441), .B2(U99_DATA1_72), 
        .ZN(n4833) );
  INV_X1 U1697 ( .A(n4832), .ZN(n4099) );
  AOI22_X1 U1698 ( .A1(n5437), .A2(n[3068]), .B1(n4733), .B2(U99_DATA1_71), 
        .ZN(n4832) );
  INV_X1 U1699 ( .A(n4831), .ZN(n4100) );
  AOI22_X1 U1700 ( .A1(n5437), .A2(n[3067]), .B1(n5438), .B2(U99_DATA1_70), 
        .ZN(n4831) );
  INV_X1 U1701 ( .A(n4830), .ZN(n4101) );
  AOI22_X1 U1702 ( .A1(n5437), .A2(n[3066]), .B1(n5439), .B2(U99_DATA1_69), 
        .ZN(n4830) );
  INV_X1 U1703 ( .A(n4829), .ZN(n4102) );
  AOI22_X1 U1704 ( .A1(n5437), .A2(n[3065]), .B1(n5440), .B2(U99_DATA1_68), 
        .ZN(n4829) );
  INV_X1 U1705 ( .A(n4828), .ZN(n4103) );
  AOI22_X1 U1706 ( .A1(n5436), .A2(n[3064]), .B1(n5440), .B2(U99_DATA1_67), 
        .ZN(n4828) );
  INV_X1 U1707 ( .A(n4827), .ZN(n4104) );
  AOI22_X1 U1708 ( .A1(n5436), .A2(n[3063]), .B1(n5440), .B2(U99_DATA1_66), 
        .ZN(n4827) );
  INV_X1 U1709 ( .A(n4826), .ZN(n4105) );
  AOI22_X1 U1710 ( .A1(n5436), .A2(n[3062]), .B1(n5440), .B2(U99_DATA1_65), 
        .ZN(n4826) );
  INV_X1 U1711 ( .A(n4825), .ZN(n4106) );
  AOI22_X1 U1712 ( .A1(n5436), .A2(n[3061]), .B1(n5440), .B2(U99_DATA1_64), 
        .ZN(n4825) );
  INV_X1 U1713 ( .A(n4824), .ZN(n4107) );
  AOI22_X1 U1714 ( .A1(n5436), .A2(n[3060]), .B1(n5440), .B2(U99_DATA1_63), 
        .ZN(n4824) );
  INV_X1 U1715 ( .A(n4823), .ZN(n4108) );
  AOI22_X1 U1716 ( .A1(n5437), .A2(n[3059]), .B1(n5440), .B2(U99_DATA1_62), 
        .ZN(n4823) );
  INV_X1 U1717 ( .A(n4822), .ZN(n4109) );
  AOI22_X1 U1718 ( .A1(n5433), .A2(n[3058]), .B1(n5439), .B2(U99_DATA1_61), 
        .ZN(n4822) );
  INV_X1 U1719 ( .A(n4821), .ZN(n4110) );
  AOI22_X1 U1720 ( .A1(n5432), .A2(n[3057]), .B1(n5439), .B2(U99_DATA1_60), 
        .ZN(n4821) );
  INV_X1 U1721 ( .A(n4820), .ZN(n4111) );
  AOI22_X1 U1722 ( .A1(n5434), .A2(n[3056]), .B1(n5439), .B2(U99_DATA1_59), 
        .ZN(n4820) );
  INV_X1 U1723 ( .A(n4819), .ZN(n4112) );
  AOI22_X1 U1724 ( .A1(n5435), .A2(n[3055]), .B1(n5439), .B2(U99_DATA1_58), 
        .ZN(n4819) );
  INV_X1 U1725 ( .A(n4818), .ZN(n4113) );
  AOI22_X1 U1726 ( .A1(n5436), .A2(n[3054]), .B1(n5439), .B2(U99_DATA1_57), 
        .ZN(n4818) );
  INV_X1 U1727 ( .A(n4817), .ZN(n4114) );
  AOI22_X1 U1728 ( .A1(n5437), .A2(n[3053]), .B1(n5438), .B2(U99_DATA1_56), 
        .ZN(n4817) );
  INV_X1 U1729 ( .A(n4816), .ZN(n4115) );
  AOI22_X1 U1730 ( .A1(n5437), .A2(n[3052]), .B1(n5438), .B2(U99_DATA1_55), 
        .ZN(n4816) );
  INV_X1 U1731 ( .A(n4815), .ZN(n4116) );
  AOI22_X1 U1732 ( .A1(n5437), .A2(n[3051]), .B1(n5438), .B2(U99_DATA1_54), 
        .ZN(n4815) );
  INV_X1 U1733 ( .A(n4814), .ZN(n4117) );
  AOI22_X1 U1734 ( .A1(n5437), .A2(n[3050]), .B1(n5438), .B2(U99_DATA1_53), 
        .ZN(n4814) );
  INV_X1 U1735 ( .A(n4813), .ZN(n4118) );
  AOI22_X1 U1736 ( .A1(n5437), .A2(n[3049]), .B1(n5438), .B2(U99_DATA1_52), 
        .ZN(n4813) );
  INV_X1 U1737 ( .A(n4804), .ZN(n4127) );
  AOI22_X1 U1738 ( .A1(n5436), .A2(n[3040]), .B1(n5431), .B2(U99_DATA1_43), 
        .ZN(n4804) );
  INV_X1 U1739 ( .A(n4803), .ZN(n4128) );
  AOI22_X1 U1740 ( .A1(n5433), .A2(n[3039]), .B1(n5441), .B2(U99_DATA1_42), 
        .ZN(n4803) );
  INV_X1 U1741 ( .A(n4802), .ZN(n4129) );
  AOI22_X1 U1742 ( .A1(n5433), .A2(n[3038]), .B1(n5431), .B2(U99_DATA1_41), 
        .ZN(n4802) );
  INV_X1 U1743 ( .A(n4801), .ZN(n4130) );
  AOI22_X1 U1744 ( .A1(n5432), .A2(n[3037]), .B1(n5441), .B2(U99_DATA1_40), 
        .ZN(n4801) );
  INV_X1 U1745 ( .A(n4800), .ZN(n4131) );
  AOI22_X1 U1746 ( .A1(n5432), .A2(n[3036]), .B1(n5441), .B2(U99_DATA1_39), 
        .ZN(n4800) );
  INV_X1 U1747 ( .A(n4799), .ZN(n4132) );
  AOI22_X1 U1748 ( .A1(n5432), .A2(n[3035]), .B1(n4733), .B2(U99_DATA1_38), 
        .ZN(n4799) );
  INV_X1 U1749 ( .A(n4798), .ZN(n4133) );
  AOI22_X1 U1750 ( .A1(n5432), .A2(n[3034]), .B1(n4733), .B2(U99_DATA1_37), 
        .ZN(n4798) );
  INV_X1 U1751 ( .A(n4797), .ZN(n4134) );
  AOI22_X1 U1752 ( .A1(n5432), .A2(n[3033]), .B1(n4733), .B2(U99_DATA1_36), 
        .ZN(n4797) );
  INV_X1 U1753 ( .A(n4796), .ZN(n4135) );
  AOI22_X1 U1754 ( .A1(n5432), .A2(n[3032]), .B1(n5441), .B2(U99_DATA1_35), 
        .ZN(n4796) );
  INV_X1 U1755 ( .A(n4795), .ZN(n4136) );
  AOI22_X1 U1756 ( .A1(n5432), .A2(n[3031]), .B1(n5439), .B2(U99_DATA1_34), 
        .ZN(n4795) );
  INV_X1 U1757 ( .A(n4794), .ZN(n4137) );
  AOI22_X1 U1758 ( .A1(n5432), .A2(n[3030]), .B1(n5440), .B2(U99_DATA1_33), 
        .ZN(n4794) );
  INV_X1 U1759 ( .A(n4793), .ZN(n4138) );
  AOI22_X1 U1760 ( .A1(n5432), .A2(n[3029]), .B1(n5440), .B2(U99_DATA1_32), 
        .ZN(n4793) );
  INV_X1 U1761 ( .A(n4792), .ZN(n4139) );
  AOI22_X1 U1762 ( .A1(n5432), .A2(n[3028]), .B1(n5431), .B2(U99_DATA1_31), 
        .ZN(n4792) );
  INV_X1 U1763 ( .A(n4791), .ZN(n4140) );
  AOI22_X1 U1764 ( .A1(n5432), .A2(n[3027]), .B1(n5441), .B2(U99_DATA1_30), 
        .ZN(n4791) );
  INV_X1 U1765 ( .A(n4790), .ZN(n4141) );
  AOI22_X1 U1766 ( .A1(n5432), .A2(n[3026]), .B1(n5441), .B2(U99_DATA1_29), 
        .ZN(n4790) );
  INV_X1 U1767 ( .A(n4789), .ZN(n4142) );
  AOI22_X1 U1768 ( .A1(n5432), .A2(n[3025]), .B1(n5441), .B2(U99_DATA1_28), 
        .ZN(n4789) );
  INV_X1 U1769 ( .A(n4788), .ZN(n4143) );
  AOI22_X1 U1770 ( .A1(n5433), .A2(n[3024]), .B1(n5441), .B2(U99_DATA1_27), 
        .ZN(n4788) );
  INV_X1 U1771 ( .A(n4787), .ZN(n4144) );
  AOI22_X1 U1772 ( .A1(n5433), .A2(n[3023]), .B1(n5438), .B2(U99_DATA1_26), 
        .ZN(n4787) );
  INV_X1 U1773 ( .A(n4786), .ZN(n4145) );
  AOI22_X1 U1774 ( .A1(n5433), .A2(n[3022]), .B1(n5441), .B2(U99_DATA1_25), 
        .ZN(n4786) );
  INV_X1 U1775 ( .A(n4785), .ZN(n4146) );
  AOI22_X1 U1776 ( .A1(n5433), .A2(n[3021]), .B1(n5431), .B2(U99_DATA1_24), 
        .ZN(n4785) );
  INV_X1 U1777 ( .A(n4784), .ZN(n4147) );
  AOI22_X1 U1778 ( .A1(n5433), .A2(n[3020]), .B1(n5431), .B2(U99_DATA1_23), 
        .ZN(n4784) );
  INV_X1 U1779 ( .A(n4783), .ZN(n4148) );
  AOI22_X1 U1780 ( .A1(n5433), .A2(n[3019]), .B1(n5441), .B2(U99_DATA1_22), 
        .ZN(n4783) );
  INV_X1 U1781 ( .A(n4782), .ZN(n4149) );
  AOI22_X1 U1782 ( .A1(n5433), .A2(n[3018]), .B1(n5441), .B2(U99_DATA1_21), 
        .ZN(n4782) );
  INV_X1 U1783 ( .A(n4781), .ZN(n4150) );
  AOI22_X1 U1784 ( .A1(n5433), .A2(n[3017]), .B1(n5439), .B2(U99_DATA1_20), 
        .ZN(n4781) );
  INV_X1 U1785 ( .A(n4780), .ZN(n4151) );
  AOI22_X1 U1786 ( .A1(n5433), .A2(n[3016]), .B1(n5441), .B2(U99_DATA1_19), 
        .ZN(n4780) );
  INV_X1 U1787 ( .A(n4779), .ZN(n4152) );
  AOI22_X1 U1788 ( .A1(n5433), .A2(n[3015]), .B1(n5439), .B2(U99_DATA1_18), 
        .ZN(n4779) );
  INV_X1 U1789 ( .A(n4778), .ZN(n4153) );
  AOI22_X1 U1790 ( .A1(n5433), .A2(n[3014]), .B1(n5438), .B2(U99_DATA1_17), 
        .ZN(n4778) );
  INV_X1 U1791 ( .A(n4777), .ZN(n4154) );
  AOI22_X1 U1792 ( .A1(n5433), .A2(n[3013]), .B1(n5441), .B2(U99_DATA1_16), 
        .ZN(n4777) );
  INV_X1 U1793 ( .A(n4776), .ZN(n4155) );
  AOI22_X1 U1794 ( .A1(n5436), .A2(n[3012]), .B1(n5440), .B2(U99_DATA1_15), 
        .ZN(n4776) );
  INV_X1 U1795 ( .A(n4775), .ZN(n4156) );
  AOI22_X1 U1796 ( .A1(n5437), .A2(n[3011]), .B1(n5438), .B2(U99_DATA1_14), 
        .ZN(n4775) );
  INV_X1 U1797 ( .A(n4774), .ZN(n4157) );
  AOI22_X1 U1798 ( .A1(n5434), .A2(n[3010]), .B1(n5431), .B2(U99_DATA1_13), 
        .ZN(n4774) );
  INV_X1 U1799 ( .A(n4773), .ZN(n4158) );
  AOI22_X1 U1800 ( .A1(n5432), .A2(n[3009]), .B1(n5431), .B2(U99_DATA1_12), 
        .ZN(n4773) );
  INV_X1 U1801 ( .A(n4772), .ZN(n4159) );
  AOI22_X1 U1802 ( .A1(n5433), .A2(n[3008]), .B1(n5439), .B2(U99_DATA1_11), 
        .ZN(n4772) );
  INV_X1 U1803 ( .A(n4771), .ZN(n4160) );
  AOI22_X1 U1804 ( .A1(n5434), .A2(n[3007]), .B1(n5438), .B2(U99_DATA1_10), 
        .ZN(n4771) );
  INV_X1 U1805 ( .A(n4770), .ZN(n4161) );
  AOI22_X1 U1806 ( .A1(n5435), .A2(n[3006]), .B1(n5441), .B2(U99_DATA1_9), 
        .ZN(n4770) );
  INV_X1 U1807 ( .A(n4769), .ZN(n4162) );
  AOI22_X1 U1808 ( .A1(n5436), .A2(n[3005]), .B1(n5431), .B2(U99_DATA1_8), 
        .ZN(n4769) );
  INV_X1 U1809 ( .A(n4768), .ZN(n4163) );
  AOI22_X1 U1810 ( .A1(n5437), .A2(n[3004]), .B1(n5441), .B2(U99_DATA1_7), 
        .ZN(n4768) );
  INV_X1 U1811 ( .A(n4767), .ZN(n4164) );
  AOI22_X1 U1812 ( .A1(n5435), .A2(n[3003]), .B1(n5441), .B2(U99_DATA1_6), 
        .ZN(n4767) );
  INV_X1 U1813 ( .A(n4766), .ZN(n4165) );
  AOI22_X1 U1814 ( .A1(n5432), .A2(n[3002]), .B1(n5441), .B2(U99_DATA1_5), 
        .ZN(n4766) );
  INV_X1 U1815 ( .A(n4765), .ZN(n4166) );
  AOI22_X1 U1816 ( .A1(n5433), .A2(n[3001]), .B1(n5441), .B2(U99_DATA1_4), 
        .ZN(n4765) );
  INV_X1 U1817 ( .A(n4764), .ZN(n4167) );
  AOI22_X1 U1818 ( .A1(n5432), .A2(n[3000]), .B1(n5440), .B2(U99_DATA1_3), 
        .ZN(n4764) );
  INV_X1 U1819 ( .A(n4763), .ZN(n4168) );
  AOI22_X1 U1820 ( .A1(n5433), .A2(n[2999]), .B1(n5438), .B2(U99_DATA1_2), 
        .ZN(n4763) );
  INV_X1 U1821 ( .A(n4762), .ZN(n4169) );
  AOI22_X1 U1822 ( .A1(n5434), .A2(n[2998]), .B1(n5438), .B2(U99_DATA1_1), 
        .ZN(n4762) );
  INV_X1 U1823 ( .A(n4761), .ZN(n4170) );
  AOI22_X1 U1824 ( .A1(n5435), .A2(n[2997]), .B1(n5441), .B2(U99_DATA1_0), 
        .ZN(n4761) );
  INV_X1 U1825 ( .A(n4867), .ZN(n4071) );
  AOI22_X1 U1826 ( .A1(n5432), .A2(n[3124]), .B1(n5438), .B2(U99_DATA1_127), 
        .ZN(n4867) );
  OAI21_X1 U1827 ( .B1(rst), .B2(n4458), .A(n5447), .ZN(n5402) );
  OAI21_X1 U1828 ( .B1(n4329), .B2(n5449), .A(n4603), .ZN(n5147) );
  NAND2_X1 U1829 ( .A1(out_data[127]), .A2(n5443), .ZN(n4603) );
  OAI21_X1 U1830 ( .B1(n5449), .B2(n4328), .A(n4604), .ZN(n5149) );
  NAND2_X1 U1831 ( .A1(out_data[126]), .A2(n4602), .ZN(n4604) );
  OAI21_X1 U1832 ( .B1(n5449), .B2(n4327), .A(n4605), .ZN(n5151) );
  NAND2_X1 U1833 ( .A1(out_data[125]), .A2(n5445), .ZN(n4605) );
  OAI21_X1 U1834 ( .B1(n5449), .B2(n4326), .A(n4606), .ZN(n5153) );
  NAND2_X1 U1835 ( .A1(out_data[124]), .A2(n5443), .ZN(n4606) );
  OAI21_X1 U1836 ( .B1(n5448), .B2(n4325), .A(n4607), .ZN(n5155) );
  NAND2_X1 U1837 ( .A1(out_data[123]), .A2(n4602), .ZN(n4607) );
  OAI21_X1 U1838 ( .B1(n5448), .B2(n4324), .A(n4608), .ZN(n5157) );
  NAND2_X1 U1839 ( .A1(out_data[122]), .A2(n5444), .ZN(n4608) );
  OAI21_X1 U1840 ( .B1(n5448), .B2(n4323), .A(n4609), .ZN(n5159) );
  NAND2_X1 U1841 ( .A1(out_data[121]), .A2(n5448), .ZN(n4609) );
  OAI21_X1 U1842 ( .B1(n5448), .B2(n4322), .A(n4610), .ZN(n5161) );
  NAND2_X1 U1843 ( .A1(out_data[120]), .A2(n5452), .ZN(n4610) );
  OAI21_X1 U1844 ( .B1(n5448), .B2(n4321), .A(n4611), .ZN(n5163) );
  NAND2_X1 U1845 ( .A1(out_data[119]), .A2(n5443), .ZN(n4611) );
  OAI21_X1 U1846 ( .B1(n5449), .B2(n4320), .A(n4612), .ZN(n5165) );
  NAND2_X1 U1847 ( .A1(out_data[118]), .A2(n5447), .ZN(n4612) );
  OAI21_X1 U1848 ( .B1(n5449), .B2(n4319), .A(n4613), .ZN(n5167) );
  NAND2_X1 U1849 ( .A1(out_data[117]), .A2(n5443), .ZN(n4613) );
  OAI21_X1 U1850 ( .B1(n5451), .B2(n4318), .A(n4614), .ZN(n5169) );
  NAND2_X1 U1851 ( .A1(out_data[116]), .A2(n5444), .ZN(n4614) );
  OAI21_X1 U1852 ( .B1(n5449), .B2(n4317), .A(n4615), .ZN(n5171) );
  NAND2_X1 U1853 ( .A1(out_data[115]), .A2(n5446), .ZN(n4615) );
  OAI21_X1 U1854 ( .B1(n5447), .B2(n4316), .A(n4616), .ZN(n5173) );
  NAND2_X1 U1855 ( .A1(out_data[114]), .A2(n5443), .ZN(n4616) );
  OAI21_X1 U1856 ( .B1(n5449), .B2(n4315), .A(n4617), .ZN(n5175) );
  NAND2_X1 U1857 ( .A1(out_data[113]), .A2(n5444), .ZN(n4617) );
  OAI21_X1 U1858 ( .B1(n5449), .B2(n4314), .A(n4618), .ZN(n5177) );
  NAND2_X1 U1859 ( .A1(out_data[112]), .A2(n5447), .ZN(n4618) );
  OAI21_X1 U1860 ( .B1(n5451), .B2(n4313), .A(n4619), .ZN(n5179) );
  NAND2_X1 U1861 ( .A1(out_data[111]), .A2(n5452), .ZN(n4619) );
  OAI21_X1 U1862 ( .B1(n5447), .B2(n4312), .A(n4620), .ZN(n5181) );
  NAND2_X1 U1863 ( .A1(out_data[110]), .A2(n4602), .ZN(n4620) );
  OAI21_X1 U1864 ( .B1(n5447), .B2(n4311), .A(n4621), .ZN(n5183) );
  NAND2_X1 U1865 ( .A1(out_data[109]), .A2(n5446), .ZN(n4621) );
  OAI21_X1 U1866 ( .B1(n5450), .B2(n4310), .A(n4622), .ZN(n5185) );
  NAND2_X1 U1867 ( .A1(out_data[108]), .A2(n5446), .ZN(n4622) );
  OAI21_X1 U1868 ( .B1(n5449), .B2(n4309), .A(n4623), .ZN(n5187) );
  NAND2_X1 U1869 ( .A1(out_data[107]), .A2(n5446), .ZN(n4623) );
  OAI21_X1 U1870 ( .B1(n5451), .B2(n4308), .A(n4624), .ZN(n5189) );
  NAND2_X1 U1871 ( .A1(out_data[106]), .A2(n5446), .ZN(n4624) );
  OAI21_X1 U1872 ( .B1(n5448), .B2(n4307), .A(n4625), .ZN(n5191) );
  NAND2_X1 U1873 ( .A1(out_data[105]), .A2(n5448), .ZN(n4625) );
  OAI21_X1 U1874 ( .B1(n5449), .B2(n4306), .A(n4626), .ZN(n5193) );
  NAND2_X1 U1875 ( .A1(out_data[104]), .A2(n5448), .ZN(n4626) );
  OAI21_X1 U1876 ( .B1(n5447), .B2(n4305), .A(n4627), .ZN(n5195) );
  NAND2_X1 U1877 ( .A1(out_data[103]), .A2(n5451), .ZN(n4627) );
  OAI21_X1 U1878 ( .B1(n5449), .B2(n4304), .A(n4628), .ZN(n5197) );
  NAND2_X1 U1879 ( .A1(out_data[102]), .A2(n5443), .ZN(n4628) );
  OAI21_X1 U1880 ( .B1(n5449), .B2(n4303), .A(n4629), .ZN(n5199) );
  NAND2_X1 U1881 ( .A1(out_data[101]), .A2(n5447), .ZN(n4629) );
  OAI21_X1 U1882 ( .B1(n5450), .B2(n4302), .A(n4630), .ZN(n5201) );
  NAND2_X1 U1883 ( .A1(out_data[100]), .A2(n5445), .ZN(n4630) );
  OAI21_X1 U1884 ( .B1(n5448), .B2(n4301), .A(n4631), .ZN(n5203) );
  NAND2_X1 U1885 ( .A1(out_data[99]), .A2(n5443), .ZN(n4631) );
  OAI21_X1 U1886 ( .B1(n5448), .B2(n4300), .A(n4632), .ZN(n5205) );
  NAND2_X1 U1887 ( .A1(out_data[98]), .A2(n5445), .ZN(n4632) );
  OAI21_X1 U1888 ( .B1(n5448), .B2(n4299), .A(n4633), .ZN(n5207) );
  NAND2_X1 U1889 ( .A1(out_data[97]), .A2(n5445), .ZN(n4633) );
  OAI21_X1 U1890 ( .B1(n5448), .B2(n4298), .A(n4634), .ZN(n5209) );
  NAND2_X1 U1891 ( .A1(out_data[96]), .A2(n5448), .ZN(n4634) );
  OAI21_X1 U1892 ( .B1(n5448), .B2(n4297), .A(n4635), .ZN(n5211) );
  NAND2_X1 U1893 ( .A1(out_data[95]), .A2(n5444), .ZN(n4635) );
  OAI21_X1 U1894 ( .B1(n5448), .B2(n4296), .A(n4636), .ZN(n5213) );
  NAND2_X1 U1895 ( .A1(out_data[94]), .A2(n5446), .ZN(n4636) );
  OAI21_X1 U1896 ( .B1(n5448), .B2(n4295), .A(n4637), .ZN(n5215) );
  NAND2_X1 U1897 ( .A1(out_data[93]), .A2(n5447), .ZN(n4637) );
  OAI21_X1 U1898 ( .B1(n5449), .B2(n4294), .A(n4638), .ZN(n5217) );
  NAND2_X1 U1899 ( .A1(out_data[92]), .A2(n5443), .ZN(n4638) );
  OAI21_X1 U1900 ( .B1(n5448), .B2(n4293), .A(n4639), .ZN(n5219) );
  NAND2_X1 U1901 ( .A1(out_data[91]), .A2(n5447), .ZN(n4639) );
  OAI21_X1 U1902 ( .B1(n5449), .B2(n4292), .A(n4640), .ZN(n5221) );
  NAND2_X1 U1903 ( .A1(out_data[90]), .A2(n5447), .ZN(n4640) );
  OAI21_X1 U1904 ( .B1(n5449), .B2(n4291), .A(n4641), .ZN(n5223) );
  NAND2_X1 U1905 ( .A1(out_data[89]), .A2(n5447), .ZN(n4641) );
  OAI21_X1 U1906 ( .B1(n5449), .B2(n4290), .A(n4642), .ZN(n5225) );
  NAND2_X1 U1907 ( .A1(out_data[88]), .A2(n5445), .ZN(n4642) );
  OAI21_X1 U1908 ( .B1(n5449), .B2(n4289), .A(n4643), .ZN(n5227) );
  NAND2_X1 U1909 ( .A1(out_data[87]), .A2(n5446), .ZN(n4643) );
  OAI21_X1 U1910 ( .B1(n5449), .B2(n4288), .A(n4644), .ZN(n5229) );
  NAND2_X1 U1911 ( .A1(out_data[86]), .A2(n5451), .ZN(n4644) );
  OAI21_X1 U1912 ( .B1(n5446), .B2(n4287), .A(n4645), .ZN(n5231) );
  NAND2_X1 U1913 ( .A1(out_data[85]), .A2(n5447), .ZN(n4645) );
  OAI21_X1 U1914 ( .B1(n5449), .B2(n4286), .A(n4646), .ZN(n5233) );
  NAND2_X1 U1915 ( .A1(out_data[84]), .A2(n5445), .ZN(n4646) );
  OAI21_X1 U1916 ( .B1(n5451), .B2(n4285), .A(n4647), .ZN(n5235) );
  NAND2_X1 U1917 ( .A1(out_data[83]), .A2(n5443), .ZN(n4647) );
  OAI21_X1 U1918 ( .B1(n5449), .B2(n4284), .A(n4648), .ZN(n5237) );
  NAND2_X1 U1919 ( .A1(out_data[82]), .A2(n5447), .ZN(n4648) );
  OAI21_X1 U1920 ( .B1(n5446), .B2(n4283), .A(n4649), .ZN(n5239) );
  NAND2_X1 U1921 ( .A1(out_data[81]), .A2(n5445), .ZN(n4649) );
  OAI21_X1 U1922 ( .B1(n5449), .B2(n4282), .A(n4650), .ZN(n5241) );
  NAND2_X1 U1923 ( .A1(out_data[80]), .A2(n5443), .ZN(n4650) );
  OAI21_X1 U1924 ( .B1(n5449), .B2(n4281), .A(n4651), .ZN(n5243) );
  NAND2_X1 U1925 ( .A1(out_data[79]), .A2(n5452), .ZN(n4651) );
  OAI21_X1 U1926 ( .B1(n5445), .B2(n4280), .A(n4652), .ZN(n5245) );
  NAND2_X1 U1927 ( .A1(out_data[78]), .A2(n5443), .ZN(n4652) );
  OAI21_X1 U1928 ( .B1(n5449), .B2(n4279), .A(n4653), .ZN(n5247) );
  NAND2_X1 U1929 ( .A1(out_data[77]), .A2(n5447), .ZN(n4653) );
  OAI21_X1 U1930 ( .B1(n5446), .B2(n4278), .A(n4654), .ZN(n5249) );
  NAND2_X1 U1931 ( .A1(out_data[76]), .A2(n5444), .ZN(n4654) );
  OAI21_X1 U1932 ( .B1(n5444), .B2(n4277), .A(n4655), .ZN(n5251) );
  NAND2_X1 U1933 ( .A1(out_data[75]), .A2(n5447), .ZN(n4655) );
  OAI21_X1 U1934 ( .B1(n5450), .B2(n4276), .A(n4656), .ZN(n5253) );
  NAND2_X1 U1935 ( .A1(out_data[74]), .A2(n5443), .ZN(n4656) );
  OAI21_X1 U1936 ( .B1(n5450), .B2(n4275), .A(n4657), .ZN(n5255) );
  NAND2_X1 U1937 ( .A1(out_data[73]), .A2(n5445), .ZN(n4657) );
  OAI21_X1 U1938 ( .B1(n5450), .B2(n4274), .A(n4658), .ZN(n5257) );
  NAND2_X1 U1939 ( .A1(out_data[72]), .A2(n5447), .ZN(n4658) );
  OAI21_X1 U1940 ( .B1(n5450), .B2(n4273), .A(n4659), .ZN(n5259) );
  NAND2_X1 U1941 ( .A1(out_data[71]), .A2(n5444), .ZN(n4659) );
  OAI21_X1 U1942 ( .B1(n5450), .B2(n4272), .A(n4660), .ZN(n5261) );
  NAND2_X1 U1943 ( .A1(out_data[70]), .A2(n5443), .ZN(n4660) );
  OAI21_X1 U1944 ( .B1(n5450), .B2(n4271), .A(n4661), .ZN(n5263) );
  NAND2_X1 U1945 ( .A1(out_data[69]), .A2(n5447), .ZN(n4661) );
  OAI21_X1 U1946 ( .B1(n5450), .B2(n4270), .A(n4662), .ZN(n5265) );
  NAND2_X1 U1947 ( .A1(out_data[68]), .A2(n5445), .ZN(n4662) );
  OAI21_X1 U1948 ( .B1(n5450), .B2(n4269), .A(n4663), .ZN(n5267) );
  NAND2_X1 U1949 ( .A1(out_data[67]), .A2(n5444), .ZN(n4663) );
  OAI21_X1 U1950 ( .B1(n5450), .B2(n4268), .A(n4664), .ZN(n5269) );
  NAND2_X1 U1951 ( .A1(out_data[66]), .A2(n5450), .ZN(n4664) );
  OAI21_X1 U1952 ( .B1(n5450), .B2(n4267), .A(n4665), .ZN(n5271) );
  NAND2_X1 U1953 ( .A1(out_data[65]), .A2(n5444), .ZN(n4665) );
  OAI21_X1 U1954 ( .B1(n5450), .B2(n4266), .A(n4666), .ZN(n5273) );
  NAND2_X1 U1955 ( .A1(out_data[64]), .A2(n5445), .ZN(n4666) );
  OAI21_X1 U1956 ( .B1(n5450), .B2(n4265), .A(n4667), .ZN(n5275) );
  NAND2_X1 U1957 ( .A1(out_data[63]), .A2(n5444), .ZN(n4667) );
  OAI21_X1 U1958 ( .B1(n5450), .B2(n4264), .A(n4668), .ZN(n5277) );
  NAND2_X1 U1959 ( .A1(out_data[62]), .A2(n5452), .ZN(n4668) );
  OAI21_X1 U1960 ( .B1(n5451), .B2(n4263), .A(n4669), .ZN(n5279) );
  NAND2_X1 U1961 ( .A1(out_data[61]), .A2(n5447), .ZN(n4669) );
  OAI21_X1 U1962 ( .B1(n5451), .B2(n4262), .A(n4670), .ZN(n5281) );
  NAND2_X1 U1963 ( .A1(out_data[60]), .A2(n5451), .ZN(n4670) );
  OAI21_X1 U1964 ( .B1(n5451), .B2(n4261), .A(n4671), .ZN(n5283) );
  NAND2_X1 U1965 ( .A1(out_data[59]), .A2(n5443), .ZN(n4671) );
  OAI21_X1 U1966 ( .B1(n5451), .B2(n4260), .A(n4672), .ZN(n5285) );
  NAND2_X1 U1967 ( .A1(out_data[58]), .A2(n5444), .ZN(n4672) );
  OAI21_X1 U1968 ( .B1(n5451), .B2(n4259), .A(n4673), .ZN(n5287) );
  NAND2_X1 U1969 ( .A1(out_data[57]), .A2(n4602), .ZN(n4673) );
  OAI21_X1 U1970 ( .B1(n5451), .B2(n4258), .A(n4674), .ZN(n5289) );
  NAND2_X1 U1971 ( .A1(out_data[56]), .A2(n4602), .ZN(n4674) );
  OAI21_X1 U1972 ( .B1(n5451), .B2(n4257), .A(n4675), .ZN(n5291) );
  NAND2_X1 U1973 ( .A1(out_data[55]), .A2(n4602), .ZN(n4675) );
  OAI21_X1 U1974 ( .B1(n5451), .B2(n4256), .A(n4676), .ZN(n5293) );
  NAND2_X1 U1975 ( .A1(out_data[54]), .A2(n4602), .ZN(n4676) );
  OAI21_X1 U1976 ( .B1(n5451), .B2(n4255), .A(n4677), .ZN(n5295) );
  NAND2_X1 U1977 ( .A1(out_data[53]), .A2(n5448), .ZN(n4677) );
  OAI21_X1 U1978 ( .B1(n5451), .B2(n4254), .A(n4678), .ZN(n5297) );
  NAND2_X1 U1979 ( .A1(out_data[52]), .A2(n5451), .ZN(n4678) );
  OAI21_X1 U1980 ( .B1(n5451), .B2(n4253), .A(n4679), .ZN(n5299) );
  NAND2_X1 U1981 ( .A1(out_data[51]), .A2(n5443), .ZN(n4679) );
  OAI21_X1 U1982 ( .B1(n5451), .B2(n4252), .A(n4680), .ZN(n5301) );
  NAND2_X1 U1983 ( .A1(out_data[50]), .A2(n5446), .ZN(n4680) );
  OAI21_X1 U1984 ( .B1(n5451), .B2(n4251), .A(n4681), .ZN(n5303) );
  NAND2_X1 U1985 ( .A1(out_data[49]), .A2(n5450), .ZN(n4681) );
  OAI21_X1 U1986 ( .B1(n5449), .B2(n4250), .A(n4682), .ZN(n5305) );
  NAND2_X1 U1987 ( .A1(out_data[48]), .A2(n5452), .ZN(n4682) );
  OAI21_X1 U1988 ( .B1(n5449), .B2(n4249), .A(n4683), .ZN(n5307) );
  NAND2_X1 U1989 ( .A1(out_data[47]), .A2(n5450), .ZN(n4683) );
  OAI21_X1 U1990 ( .B1(n5449), .B2(n4248), .A(n4684), .ZN(n5309) );
  NAND2_X1 U1991 ( .A1(out_data[46]), .A2(n5448), .ZN(n4684) );
  OAI21_X1 U1992 ( .B1(n5449), .B2(n4247), .A(n4685), .ZN(n5311) );
  NAND2_X1 U1993 ( .A1(out_data[45]), .A2(n5446), .ZN(n4685) );
  OAI21_X1 U1994 ( .B1(n5449), .B2(n4246), .A(n4686), .ZN(n5313) );
  NAND2_X1 U1995 ( .A1(out_data[44]), .A2(n5446), .ZN(n4686) );
  OAI21_X1 U1996 ( .B1(n5452), .B2(n4245), .A(n4687), .ZN(n5315) );
  NAND2_X1 U1997 ( .A1(out_data[43]), .A2(n5446), .ZN(n4687) );
  OAI21_X1 U1998 ( .B1(n5452), .B2(n4244), .A(n4688), .ZN(n5317) );
  NAND2_X1 U1999 ( .A1(out_data[42]), .A2(n5446), .ZN(n4688) );
  OAI21_X1 U2000 ( .B1(n5452), .B2(n4243), .A(n4689), .ZN(n5319) );
  NAND2_X1 U2001 ( .A1(out_data[41]), .A2(n5446), .ZN(n4689) );
  OAI21_X1 U2002 ( .B1(n5452), .B2(n4242), .A(n4690), .ZN(n5321) );
  NAND2_X1 U2003 ( .A1(out_data[40]), .A2(n5446), .ZN(n4690) );
  OAI21_X1 U2004 ( .B1(n5452), .B2(n4241), .A(n4691), .ZN(n5323) );
  NAND2_X1 U2005 ( .A1(out_data[39]), .A2(n5446), .ZN(n4691) );
  OAI21_X1 U2006 ( .B1(n5452), .B2(n4240), .A(n4692), .ZN(n5325) );
  NAND2_X1 U2007 ( .A1(out_data[38]), .A2(n5446), .ZN(n4692) );
  OAI21_X1 U2008 ( .B1(n5452), .B2(n4239), .A(n4693), .ZN(n5327) );
  NAND2_X1 U2009 ( .A1(out_data[37]), .A2(n5446), .ZN(n4693) );
  OAI21_X1 U2010 ( .B1(n5452), .B2(n4238), .A(n4694), .ZN(n5329) );
  NAND2_X1 U2011 ( .A1(out_data[36]), .A2(n5448), .ZN(n4694) );
  OAI21_X1 U2012 ( .B1(n5445), .B2(n4237), .A(n4695), .ZN(n5331) );
  NAND2_X1 U2013 ( .A1(out_data[35]), .A2(n5446), .ZN(n4695) );
  OAI21_X1 U2014 ( .B1(n5452), .B2(n4236), .A(n4696), .ZN(n5333) );
  NAND2_X1 U2015 ( .A1(out_data[34]), .A2(n5443), .ZN(n4696) );
  OAI21_X1 U2016 ( .B1(n5449), .B2(n4235), .A(n4697), .ZN(n5335) );
  NAND2_X1 U2017 ( .A1(out_data[33]), .A2(n5447), .ZN(n4697) );
  OAI21_X1 U2018 ( .B1(n5445), .B2(n4234), .A(n4698), .ZN(n5337) );
  NAND2_X1 U2019 ( .A1(out_data[32]), .A2(n5451), .ZN(n4698) );
  OAI21_X1 U2020 ( .B1(n5448), .B2(n4233), .A(n4699), .ZN(n5339) );
  NAND2_X1 U2021 ( .A1(out_data[31]), .A2(n5447), .ZN(n4699) );
  OAI21_X1 U2022 ( .B1(n5444), .B2(n4232), .A(n4700), .ZN(n5341) );
  NAND2_X1 U2023 ( .A1(out_data[30]), .A2(n5447), .ZN(n4700) );
  OAI21_X1 U2024 ( .B1(n5450), .B2(n4231), .A(n4701), .ZN(n5343) );
  NAND2_X1 U2025 ( .A1(out_data[29]), .A2(n5443), .ZN(n4701) );
  OAI21_X1 U2026 ( .B1(n5450), .B2(n4230), .A(n4702), .ZN(n5345) );
  NAND2_X1 U2027 ( .A1(out_data[28]), .A2(n5447), .ZN(n4702) );
  OAI21_X1 U2028 ( .B1(n5447), .B2(n4229), .A(n4703), .ZN(n5347) );
  NAND2_X1 U2029 ( .A1(out_data[27]), .A2(n4602), .ZN(n4703) );
  OAI21_X1 U2030 ( .B1(n5446), .B2(n4228), .A(n4704), .ZN(n5349) );
  NAND2_X1 U2031 ( .A1(out_data[26]), .A2(n5443), .ZN(n4704) );
  OAI21_X1 U2032 ( .B1(n5447), .B2(n4227), .A(n4705), .ZN(n5351) );
  NAND2_X1 U2033 ( .A1(out_data[25]), .A2(n5443), .ZN(n4705) );
  OAI21_X1 U2034 ( .B1(n5445), .B2(n4226), .A(n4706), .ZN(n5353) );
  NAND2_X1 U2035 ( .A1(out_data[24]), .A2(n4602), .ZN(n4706) );
  OAI21_X1 U2036 ( .B1(n5447), .B2(n4225), .A(n4707), .ZN(n5355) );
  NAND2_X1 U2037 ( .A1(out_data[23]), .A2(n5447), .ZN(n4707) );
  OAI21_X1 U2038 ( .B1(n5444), .B2(n4224), .A(n4708), .ZN(n5357) );
  NAND2_X1 U2039 ( .A1(out_data[22]), .A2(n5444), .ZN(n4708) );
  OAI21_X1 U2040 ( .B1(n4602), .B2(n4223), .A(n4709), .ZN(n5359) );
  NAND2_X1 U2041 ( .A1(out_data[21]), .A2(n4602), .ZN(n4709) );
  OAI21_X1 U2042 ( .B1(n4602), .B2(n4222), .A(n4710), .ZN(n5361) );
  NAND2_X1 U2043 ( .A1(out_data[20]), .A2(n5451), .ZN(n4710) );
  OAI21_X1 U2044 ( .B1(n4602), .B2(n4221), .A(n4711), .ZN(n5363) );
  NAND2_X1 U2045 ( .A1(out_data[19]), .A2(n4602), .ZN(n4711) );
  OAI21_X1 U2046 ( .B1(n4602), .B2(n4220), .A(n4712), .ZN(n5365) );
  NAND2_X1 U2047 ( .A1(out_data[18]), .A2(n5443), .ZN(n4712) );
  OAI21_X1 U2048 ( .B1(n5450), .B2(n4219), .A(n4713), .ZN(n5367) );
  NAND2_X1 U2049 ( .A1(out_data[17]), .A2(n5443), .ZN(n4713) );
  OAI21_X1 U2050 ( .B1(n5452), .B2(n4218), .A(n4714), .ZN(n5369) );
  NAND2_X1 U2051 ( .A1(out_data[16]), .A2(n5451), .ZN(n4714) );
  OAI21_X1 U2052 ( .B1(n4602), .B2(n4217), .A(n4715), .ZN(n5371) );
  NAND2_X1 U2053 ( .A1(out_data[15]), .A2(n5445), .ZN(n4715) );
  OAI21_X1 U2054 ( .B1(n5447), .B2(n4216), .A(n4716), .ZN(n5373) );
  NAND2_X1 U2055 ( .A1(out_data[14]), .A2(n5445), .ZN(n4716) );
  OAI21_X1 U2056 ( .B1(n4602), .B2(n4215), .A(n4717), .ZN(n5375) );
  NAND2_X1 U2057 ( .A1(out_data[13]), .A2(n5445), .ZN(n4717) );
  OAI21_X1 U2058 ( .B1(n4602), .B2(n4214), .A(n4718), .ZN(n5377) );
  NAND2_X1 U2059 ( .A1(out_data[12]), .A2(n5447), .ZN(n4718) );
  OAI21_X1 U2060 ( .B1(n5444), .B2(n4213), .A(n4719), .ZN(n5379) );
  NAND2_X1 U2061 ( .A1(out_data[11]), .A2(n5447), .ZN(n4719) );
  OAI21_X1 U2062 ( .B1(n5448), .B2(n4212), .A(n4720), .ZN(n5381) );
  NAND2_X1 U2063 ( .A1(out_data[10]), .A2(n5446), .ZN(n4720) );
  OAI21_X1 U2064 ( .B1(n5452), .B2(n4211), .A(n4721), .ZN(n5383) );
  NAND2_X1 U2065 ( .A1(out_data[9]), .A2(n5447), .ZN(n4721) );
  OAI21_X1 U2066 ( .B1(n5448), .B2(n4210), .A(n4722), .ZN(n5385) );
  NAND2_X1 U2067 ( .A1(out_data[8]), .A2(n5444), .ZN(n4722) );
  OAI21_X1 U2068 ( .B1(n5445), .B2(n4209), .A(n4723), .ZN(n5387) );
  NAND2_X1 U2069 ( .A1(out_data[7]), .A2(n5451), .ZN(n4723) );
  OAI21_X1 U2070 ( .B1(n5444), .B2(n4208), .A(n4724), .ZN(n5389) );
  NAND2_X1 U2071 ( .A1(out_data[6]), .A2(n5443), .ZN(n4724) );
  OAI21_X1 U2072 ( .B1(n5450), .B2(n4207), .A(n4725), .ZN(n5391) );
  NAND2_X1 U2073 ( .A1(out_data[5]), .A2(n5444), .ZN(n4725) );
  OAI21_X1 U2074 ( .B1(n5449), .B2(n4206), .A(n4726), .ZN(n5393) );
  NAND2_X1 U2075 ( .A1(out_data[4]), .A2(n5444), .ZN(n4726) );
  OAI21_X1 U2076 ( .B1(n5444), .B2(n4205), .A(n4727), .ZN(n5395) );
  NAND2_X1 U2077 ( .A1(out_data[3]), .A2(n5450), .ZN(n4727) );
  OAI21_X1 U2078 ( .B1(n5445), .B2(n4204), .A(n4728), .ZN(n5397) );
  NAND2_X1 U2079 ( .A1(out_data[2]), .A2(n5445), .ZN(n4728) );
  OAI21_X1 U2080 ( .B1(n4602), .B2(n4203), .A(n4729), .ZN(n5399) );
  NAND2_X1 U2081 ( .A1(out_data[1]), .A2(n5444), .ZN(n4729) );
  OAI21_X1 U2082 ( .B1(n5449), .B2(n4202), .A(n4731), .ZN(n5401) );
  NAND2_X1 U2083 ( .A1(out_data[0]), .A2(n5445), .ZN(n4731) );
  INV_X1 U2084 ( .A(rst), .ZN(n4600) );
  INV_X1 U2085 ( .A(n3389), .ZN(n4328) );
  INV_X1 U2086 ( .A(n3388), .ZN(n4327) );
  INV_X1 U2087 ( .A(n3387), .ZN(n4326) );
  INV_X1 U2088 ( .A(n3386), .ZN(n4325) );
  INV_X1 U2089 ( .A(n3385), .ZN(n4324) );
  INV_X1 U2090 ( .A(n3384), .ZN(n4323) );
  INV_X1 U2091 ( .A(n3383), .ZN(n4322) );
  INV_X1 U2092 ( .A(n3382), .ZN(n4321) );
  INV_X1 U2093 ( .A(n3381), .ZN(n4320) );
  INV_X1 U2094 ( .A(n3380), .ZN(n4319) );
  INV_X1 U2095 ( .A(n3379), .ZN(n4318) );
  INV_X1 U2096 ( .A(n3378), .ZN(n4317) );
  INV_X1 U2097 ( .A(n3377), .ZN(n4316) );
  INV_X1 U2098 ( .A(n3376), .ZN(n4315) );
  INV_X1 U2099 ( .A(n3375), .ZN(n4314) );
  INV_X1 U2100 ( .A(n3374), .ZN(n4313) );
  INV_X1 U2101 ( .A(n3373), .ZN(n4312) );
  INV_X1 U2102 ( .A(n3372), .ZN(n4311) );
  INV_X1 U2103 ( .A(n3371), .ZN(n4310) );
  INV_X1 U2104 ( .A(n3370), .ZN(n4309) );
  INV_X1 U2105 ( .A(n3369), .ZN(n4308) );
  INV_X1 U2106 ( .A(n3368), .ZN(n4307) );
  INV_X1 U2107 ( .A(n3367), .ZN(n4306) );
  INV_X1 U2108 ( .A(n3366), .ZN(n4305) );
  INV_X1 U2109 ( .A(n3365), .ZN(n4304) );
  INV_X1 U2110 ( .A(n3364), .ZN(n4303) );
  INV_X1 U2111 ( .A(n3363), .ZN(n4302) );
  INV_X1 U2112 ( .A(n3362), .ZN(n4301) );
  INV_X1 U2113 ( .A(n3361), .ZN(n4300) );
  INV_X1 U2114 ( .A(n3360), .ZN(n4299) );
  INV_X1 U2115 ( .A(n3359), .ZN(n4298) );
  INV_X1 U2116 ( .A(n3358), .ZN(n4297) );
  INV_X1 U2117 ( .A(n3357), .ZN(n4296) );
  INV_X1 U2118 ( .A(n3356), .ZN(n4295) );
  INV_X1 U2119 ( .A(n3355), .ZN(n4294) );
  INV_X1 U2120 ( .A(n3354), .ZN(n4293) );
  INV_X1 U2121 ( .A(n3353), .ZN(n4292) );
  INV_X1 U2122 ( .A(n3352), .ZN(n4291) );
  INV_X1 U2123 ( .A(n3351), .ZN(n4290) );
  INV_X1 U2124 ( .A(n3350), .ZN(n4289) );
  INV_X1 U2125 ( .A(n3349), .ZN(n4288) );
  INV_X1 U2126 ( .A(n3348), .ZN(n4287) );
  INV_X1 U2127 ( .A(n3347), .ZN(n4286) );
  INV_X1 U2128 ( .A(n3346), .ZN(n4285) );
  INV_X1 U2129 ( .A(n3345), .ZN(n4284) );
  INV_X1 U2130 ( .A(n3344), .ZN(n4283) );
  INV_X1 U2131 ( .A(n3343), .ZN(n4282) );
  INV_X1 U2132 ( .A(n3342), .ZN(n4281) );
  INV_X1 U2133 ( .A(n3341), .ZN(n4280) );
  INV_X1 U2134 ( .A(n3340), .ZN(n4279) );
  INV_X1 U2135 ( .A(n3339), .ZN(n4278) );
  INV_X1 U2136 ( .A(n3338), .ZN(n4277) );
  INV_X1 U2137 ( .A(n3337), .ZN(n4276) );
  INV_X1 U2138 ( .A(n3336), .ZN(n4275) );
  INV_X1 U2139 ( .A(n3335), .ZN(n4274) );
  INV_X1 U2140 ( .A(n3334), .ZN(n4273) );
  INV_X1 U2141 ( .A(n3333), .ZN(n4272) );
  INV_X1 U2142 ( .A(n3332), .ZN(n4271) );
  INV_X1 U2143 ( .A(n3331), .ZN(n4270) );
  INV_X1 U2144 ( .A(n3330), .ZN(n4269) );
  INV_X1 U2145 ( .A(n3329), .ZN(n4268) );
  INV_X1 U2146 ( .A(n3328), .ZN(n4267) );
  INV_X1 U2147 ( .A(n3327), .ZN(n4266) );
  INV_X1 U2148 ( .A(n3326), .ZN(n4265) );
  INV_X1 U2149 ( .A(n3325), .ZN(n4264) );
  INV_X1 U2150 ( .A(n3324), .ZN(n4263) );
  INV_X1 U2151 ( .A(n3323), .ZN(n4262) );
  INV_X1 U2152 ( .A(n3322), .ZN(n4261) );
  INV_X1 U2153 ( .A(n3321), .ZN(n4260) );
  INV_X1 U2154 ( .A(n3320), .ZN(n4259) );
  INV_X1 U2155 ( .A(n3319), .ZN(n4258) );
  INV_X1 U2156 ( .A(n3318), .ZN(n4257) );
  INV_X1 U2157 ( .A(n3317), .ZN(n4256) );
  INV_X1 U2158 ( .A(n3316), .ZN(n4255) );
  INV_X1 U2159 ( .A(n3315), .ZN(n4254) );
  INV_X1 U2160 ( .A(n3314), .ZN(n4253) );
  INV_X1 U2161 ( .A(n3313), .ZN(n4252) );
  INV_X1 U2162 ( .A(n3312), .ZN(n4251) );
  INV_X1 U2163 ( .A(n3311), .ZN(n4250) );
  INV_X1 U2164 ( .A(n3310), .ZN(n4249) );
  INV_X1 U2165 ( .A(n3309), .ZN(n4248) );
  INV_X1 U2166 ( .A(n3308), .ZN(n4247) );
  INV_X1 U2167 ( .A(n3307), .ZN(n4246) );
  INV_X1 U2168 ( .A(n3306), .ZN(n4245) );
  INV_X1 U2169 ( .A(n3305), .ZN(n4244) );
  INV_X1 U2170 ( .A(n3304), .ZN(n4243) );
  INV_X1 U2171 ( .A(n3303), .ZN(n4242) );
  INV_X1 U2172 ( .A(n3302), .ZN(n4241) );
  INV_X1 U2173 ( .A(n3301), .ZN(n4240) );
  INV_X1 U2174 ( .A(n3300), .ZN(n4239) );
  INV_X1 U2175 ( .A(n3299), .ZN(n4238) );
  INV_X1 U2176 ( .A(n3298), .ZN(n4237) );
  INV_X1 U2177 ( .A(n3297), .ZN(n4236) );
  INV_X1 U2178 ( .A(n3296), .ZN(n4235) );
  INV_X1 U2179 ( .A(n3295), .ZN(n4234) );
  INV_X1 U2180 ( .A(n3294), .ZN(n4233) );
  INV_X1 U2181 ( .A(n3293), .ZN(n4232) );
  INV_X1 U2182 ( .A(n3292), .ZN(n4231) );
  INV_X1 U2183 ( .A(n3291), .ZN(n4230) );
  INV_X1 U2184 ( .A(n3290), .ZN(n4229) );
  INV_X1 U2185 ( .A(n3289), .ZN(n4228) );
  INV_X1 U2186 ( .A(n3288), .ZN(n4227) );
  INV_X1 U2187 ( .A(n3287), .ZN(n4226) );
  INV_X1 U2188 ( .A(n3286), .ZN(n4225) );
  INV_X1 U2189 ( .A(n3285), .ZN(n4224) );
  INV_X1 U2190 ( .A(n3284), .ZN(n4223) );
  INV_X1 U2191 ( .A(n3283), .ZN(n4222) );
  INV_X1 U2192 ( .A(n3282), .ZN(n4221) );
  INV_X1 U2193 ( .A(n3281), .ZN(n4220) );
  INV_X1 U2194 ( .A(n3280), .ZN(n4219) );
  INV_X1 U2195 ( .A(n3279), .ZN(n4218) );
  INV_X1 U2196 ( .A(n3278), .ZN(n4217) );
  INV_X1 U2197 ( .A(n3277), .ZN(n4216) );
  INV_X1 U2198 ( .A(n3276), .ZN(n4215) );
  INV_X1 U2199 ( .A(n3275), .ZN(n4214) );
  INV_X1 U2200 ( .A(n3274), .ZN(n4213) );
  INV_X1 U2201 ( .A(n3273), .ZN(n4212) );
  INV_X1 U2202 ( .A(n3272), .ZN(n4211) );
  INV_X1 U2203 ( .A(n3271), .ZN(n4210) );
  INV_X1 U2204 ( .A(n3270), .ZN(n4209) );
  INV_X1 U2205 ( .A(n3269), .ZN(n4208) );
  INV_X1 U2206 ( .A(n3268), .ZN(n4207) );
  INV_X1 U2207 ( .A(n3267), .ZN(n4206) );
  INV_X1 U2208 ( .A(n3266), .ZN(n4205) );
  INV_X1 U2209 ( .A(n3265), .ZN(n4204) );
  INV_X1 U2210 ( .A(n3264), .ZN(n4203) );
  INV_X1 U2211 ( .A(n3263), .ZN(n4202) );
  INV_X1 U2212 ( .A(n3390), .ZN(n4329) );
  OAI22_X1 U2214 ( .A1(n5415), .A2(n4462), .B1(n5107), .B2(n5410), .ZN(
        U49_Z_127) );
  XNOR2_X1 U2215 ( .A(key_in[127]), .B(data_in[127]), .ZN(n5107) );
  OAI22_X1 U2216 ( .A1(n5415), .A2(n4463), .B1(n5108), .B2(n5413), .ZN(
        U49_Z_126) );
  XNOR2_X1 U2217 ( .A(key_in[126]), .B(data_in[126]), .ZN(n5108) );
  OAI22_X1 U2218 ( .A1(n5415), .A2(n4464), .B1(n5109), .B2(n5412), .ZN(
        U49_Z_125) );
  XNOR2_X1 U2219 ( .A(key_in[125]), .B(data_in[125]), .ZN(n5109) );
  OAI22_X1 U2220 ( .A1(n5419), .A2(n4465), .B1(n5110), .B2(n5413), .ZN(
        U49_Z_124) );
  XNOR2_X1 U2221 ( .A(key_in[124]), .B(data_in[124]), .ZN(n5110) );
  OAI22_X1 U2222 ( .A1(n5416), .A2(n4466), .B1(n5111), .B2(n5409), .ZN(
        U49_Z_123) );
  XNOR2_X1 U2223 ( .A(key_in[123]), .B(data_in[123]), .ZN(n5111) );
  OAI22_X1 U2224 ( .A1(n5418), .A2(n4467), .B1(n5112), .B2(n5412), .ZN(
        U49_Z_122) );
  XNOR2_X1 U2225 ( .A(key_in[122]), .B(data_in[122]), .ZN(n5112) );
  OAI22_X1 U2226 ( .A1(n5416), .A2(n4566), .B1(n5095), .B2(n5412), .ZN(
        U49_Z_23) );
  XNOR2_X1 U2227 ( .A(key_in[23]), .B(data_in[23]), .ZN(n5095) );
  OAI22_X1 U2228 ( .A1(n5416), .A2(n4567), .B1(n5096), .B2(n5413), .ZN(
        U49_Z_22) );
  XNOR2_X1 U2229 ( .A(key_in[22]), .B(data_in[22]), .ZN(n5096) );
  OAI22_X1 U2230 ( .A1(n5416), .A2(n4568), .B1(n5097), .B2(n5412), .ZN(
        U49_Z_21) );
  XNOR2_X1 U2231 ( .A(key_in[21]), .B(data_in[21]), .ZN(n5097) );
  OAI22_X1 U2232 ( .A1(n5416), .A2(n4569), .B1(n5098), .B2(n5410), .ZN(
        U49_Z_20) );
  XNOR2_X1 U2233 ( .A(key_in[20]), .B(data_in[20]), .ZN(n5098) );
  OAI22_X1 U2234 ( .A1(n5415), .A2(n4570), .B1(n5100), .B2(n5409), .ZN(
        U49_Z_19) );
  XNOR2_X1 U2235 ( .A(key_in[19]), .B(data_in[19]), .ZN(n5100) );
  OAI22_X1 U2236 ( .A1(n5415), .A2(n4571), .B1(n5101), .B2(n5411), .ZN(
        U49_Z_18) );
  XNOR2_X1 U2237 ( .A(key_in[18]), .B(data_in[18]), .ZN(n5101) );
  OAI22_X1 U2238 ( .A1(n5416), .A2(n4572), .B1(n5102), .B2(n5412), .ZN(
        U49_Z_17) );
  XNOR2_X1 U2239 ( .A(key_in[17]), .B(data_in[17]), .ZN(n5102) );
  OAI22_X1 U2240 ( .A1(n5417), .A2(n4573), .B1(n5103), .B2(n5413), .ZN(
        U49_Z_16) );
  XNOR2_X1 U2241 ( .A(key_in[16]), .B(data_in[16]), .ZN(n5103) );
  OAI22_X1 U2242 ( .A1(n5418), .A2(n4574), .B1(n5104), .B2(n5413), .ZN(
        U49_Z_15) );
  XNOR2_X1 U2243 ( .A(key_in[15]), .B(data_in[15]), .ZN(n5104) );
  OAI22_X1 U2244 ( .A1(n5415), .A2(n4575), .B1(n5105), .B2(n5411), .ZN(
        U49_Z_14) );
  XNOR2_X1 U2245 ( .A(key_in[14]), .B(data_in[14]), .ZN(n5105) );
  OAI22_X1 U2246 ( .A1(n5415), .A2(n4576), .B1(n5106), .B2(n5409), .ZN(
        U49_Z_13) );
  XNOR2_X1 U2247 ( .A(key_in[13]), .B(data_in[13]), .ZN(n5106) );
  OAI22_X1 U2248 ( .A1(n5416), .A2(n4587), .B1(n5099), .B2(n5411), .ZN(U49_Z_2) );
  XNOR2_X1 U2249 ( .A(key_in[2]), .B(data_in[2]), .ZN(n5099) );
  AOI21_X1 U2250 ( .B1(n5142), .B2(n5143), .A(ready), .ZN(U47_Z_1) );
  OAI22_X1 U2251 ( .A1(n5415), .A2(n4490), .B1(n5011), .B2(n5012), .ZN(
        U49_Z_99) );
  XNOR2_X1 U2252 ( .A(key_in[99]), .B(data_in[99]), .ZN(n5011) );
  OAI22_X1 U2253 ( .A1(n5419), .A2(n4491), .B1(n5013), .B2(n5012), .ZN(
        U49_Z_98) );
  XNOR2_X1 U2254 ( .A(key_in[98]), .B(data_in[98]), .ZN(n5013) );
  OAI22_X1 U2255 ( .A1(n5419), .A2(n4492), .B1(n5014), .B2(n5413), .ZN(
        U49_Z_97) );
  XNOR2_X1 U2256 ( .A(key_in[97]), .B(data_in[97]), .ZN(n5014) );
  OAI22_X1 U2257 ( .A1(n5418), .A2(n4493), .B1(n5015), .B2(n5413), .ZN(
        U49_Z_96) );
  XNOR2_X1 U2258 ( .A(key_in[96]), .B(data_in[96]), .ZN(n5015) );
  OAI22_X1 U2259 ( .A1(n5418), .A2(n4494), .B1(n5016), .B2(n5413), .ZN(
        U49_Z_95) );
  XNOR2_X1 U2260 ( .A(key_in[95]), .B(data_in[95]), .ZN(n5016) );
  OAI22_X1 U2261 ( .A1(n5418), .A2(n4495), .B1(n5017), .B2(n5413), .ZN(
        U49_Z_94) );
  XNOR2_X1 U2262 ( .A(key_in[94]), .B(data_in[94]), .ZN(n5017) );
  OAI22_X1 U2263 ( .A1(n5418), .A2(n4496), .B1(n5018), .B2(n5413), .ZN(
        U49_Z_93) );
  XNOR2_X1 U2264 ( .A(key_in[93]), .B(data_in[93]), .ZN(n5018) );
  OAI22_X1 U2265 ( .A1(n5418), .A2(n4497), .B1(n5019), .B2(n5413), .ZN(
        U49_Z_92) );
  XNOR2_X1 U2266 ( .A(key_in[92]), .B(data_in[92]), .ZN(n5019) );
  OAI22_X1 U2267 ( .A1(n5418), .A2(n4498), .B1(n5020), .B2(n5413), .ZN(
        U49_Z_91) );
  XNOR2_X1 U2268 ( .A(key_in[91]), .B(data_in[91]), .ZN(n5020) );
  OAI22_X1 U2269 ( .A1(n5417), .A2(n4499), .B1(n5021), .B2(n5413), .ZN(
        U49_Z_90) );
  XNOR2_X1 U2270 ( .A(key_in[90]), .B(data_in[90]), .ZN(n5021) );
  OAI22_X1 U2271 ( .A1(n5415), .A2(n4500), .B1(n5023), .B2(n5412), .ZN(
        U49_Z_89) );
  XNOR2_X1 U2272 ( .A(key_in[89]), .B(data_in[89]), .ZN(n5023) );
  OAI22_X1 U2273 ( .A1(n5417), .A2(n4501), .B1(n5024), .B2(n5412), .ZN(
        U49_Z_88) );
  XNOR2_X1 U2274 ( .A(key_in[88]), .B(data_in[88]), .ZN(n5024) );
  OAI22_X1 U2275 ( .A1(n5418), .A2(n4502), .B1(n5025), .B2(n5412), .ZN(
        U49_Z_87) );
  XNOR2_X1 U2276 ( .A(key_in[87]), .B(data_in[87]), .ZN(n5025) );
  OAI22_X1 U2277 ( .A1(n5418), .A2(n4503), .B1(n5026), .B2(n5412), .ZN(
        U49_Z_86) );
  XNOR2_X1 U2278 ( .A(key_in[86]), .B(data_in[86]), .ZN(n5026) );
  OAI22_X1 U2279 ( .A1(n5416), .A2(n4504), .B1(n5027), .B2(n5412), .ZN(
        U49_Z_85) );
  XNOR2_X1 U2280 ( .A(key_in[85]), .B(data_in[85]), .ZN(n5027) );
  OAI22_X1 U2281 ( .A1(n5417), .A2(n4505), .B1(n5028), .B2(n5412), .ZN(
        U49_Z_84) );
  XNOR2_X1 U2282 ( .A(key_in[84]), .B(data_in[84]), .ZN(n5028) );
  OAI22_X1 U2283 ( .A1(n5416), .A2(n4506), .B1(n5029), .B2(n5412), .ZN(
        U49_Z_83) );
  XNOR2_X1 U2284 ( .A(key_in[83]), .B(data_in[83]), .ZN(n5029) );
  OAI22_X1 U2285 ( .A1(n5419), .A2(n4507), .B1(n5030), .B2(n5412), .ZN(
        U49_Z_82) );
  XNOR2_X1 U2286 ( .A(key_in[82]), .B(data_in[82]), .ZN(n5030) );
  OAI22_X1 U2287 ( .A1(n5416), .A2(n4508), .B1(n5031), .B2(n5412), .ZN(
        U49_Z_81) );
  XNOR2_X1 U2288 ( .A(key_in[81]), .B(data_in[81]), .ZN(n5031) );
  OAI22_X1 U2289 ( .A1(n5417), .A2(n4509), .B1(n5032), .B2(n5411), .ZN(
        U49_Z_80) );
  XNOR2_X1 U2290 ( .A(key_in[80]), .B(data_in[80]), .ZN(n5032) );
  OAI22_X1 U2291 ( .A1(n5416), .A2(n4510), .B1(n5034), .B2(n5411), .ZN(
        U49_Z_79) );
  XNOR2_X1 U2292 ( .A(key_in[79]), .B(data_in[79]), .ZN(n5034) );
  OAI22_X1 U2293 ( .A1(n5417), .A2(n4511), .B1(n5035), .B2(n5411), .ZN(
        U49_Z_78) );
  XNOR2_X1 U2294 ( .A(key_in[78]), .B(data_in[78]), .ZN(n5035) );
  OAI22_X1 U2295 ( .A1(n5419), .A2(n4512), .B1(n5036), .B2(n5411), .ZN(
        U49_Z_77) );
  XNOR2_X1 U2296 ( .A(key_in[77]), .B(data_in[77]), .ZN(n5036) );
  OAI22_X1 U2297 ( .A1(n5415), .A2(n4513), .B1(n5037), .B2(n5411), .ZN(
        U49_Z_76) );
  XNOR2_X1 U2298 ( .A(key_in[76]), .B(data_in[76]), .ZN(n5037) );
  OAI22_X1 U2299 ( .A1(n5414), .A2(n4514), .B1(n5038), .B2(n5411), .ZN(
        U49_Z_75) );
  XNOR2_X1 U2300 ( .A(key_in[75]), .B(data_in[75]), .ZN(n5038) );
  OAI22_X1 U2301 ( .A1(n5419), .A2(n4515), .B1(n5039), .B2(n5411), .ZN(
        U49_Z_74) );
  XNOR2_X1 U2302 ( .A(key_in[74]), .B(data_in[74]), .ZN(n5039) );
  OAI22_X1 U2303 ( .A1(n5414), .A2(n4516), .B1(n5040), .B2(n5411), .ZN(
        U49_Z_73) );
  XNOR2_X1 U2304 ( .A(key_in[73]), .B(data_in[73]), .ZN(n5040) );
  OAI22_X1 U2305 ( .A1(n5415), .A2(n4580), .B1(n5022), .B2(n5413), .ZN(U49_Z_9) );
  XNOR2_X1 U2306 ( .A(key_in[9]), .B(data_in[9]), .ZN(n5022) );
  OAI22_X1 U2307 ( .A1(n5414), .A2(n4581), .B1(n5033), .B2(n5411), .ZN(U49_Z_8) );
  XNOR2_X1 U2308 ( .A(key_in[8]), .B(data_in[8]), .ZN(n5033) );
  OAI22_X1 U2309 ( .A1(n5419), .A2(n4468), .B1(n5113), .B2(n5410), .ZN(
        U49_Z_121) );
  XNOR2_X1 U2310 ( .A(key_in[121]), .B(data_in[121]), .ZN(n5113) );
  OAI22_X1 U2311 ( .A1(n5418), .A2(n4469), .B1(n5114), .B2(n5410), .ZN(
        U49_Z_120) );
  XNOR2_X1 U2312 ( .A(key_in[120]), .B(data_in[120]), .ZN(n5114) );
  OAI22_X1 U2313 ( .A1(n5414), .A2(n4470), .B1(n5116), .B2(n5410), .ZN(
        U49_Z_119) );
  XNOR2_X1 U2314 ( .A(key_in[119]), .B(data_in[119]), .ZN(n5116) );
  OAI22_X1 U2315 ( .A1(n5414), .A2(n4471), .B1(n5117), .B2(n5410), .ZN(
        U49_Z_118) );
  XNOR2_X1 U2316 ( .A(key_in[118]), .B(data_in[118]), .ZN(n5117) );
  OAI22_X1 U2317 ( .A1(n5414), .A2(n4472), .B1(n5118), .B2(n5410), .ZN(
        U49_Z_117) );
  XNOR2_X1 U2318 ( .A(key_in[117]), .B(data_in[117]), .ZN(n5118) );
  OAI22_X1 U2319 ( .A1(n5414), .A2(n4473), .B1(n5119), .B2(n5410), .ZN(
        U49_Z_116) );
  XNOR2_X1 U2320 ( .A(key_in[116]), .B(data_in[116]), .ZN(n5119) );
  OAI22_X1 U2321 ( .A1(n5416), .A2(n4474), .B1(n5120), .B2(n5410), .ZN(
        U49_Z_115) );
  XNOR2_X1 U2322 ( .A(key_in[115]), .B(data_in[115]), .ZN(n5120) );
  OAI22_X1 U2323 ( .A1(n5416), .A2(n4475), .B1(n5121), .B2(n5410), .ZN(
        U49_Z_114) );
  XNOR2_X1 U2324 ( .A(key_in[114]), .B(data_in[114]), .ZN(n5121) );
  OAI22_X1 U2325 ( .A1(n5415), .A2(n4476), .B1(n5122), .B2(n5409), .ZN(
        U49_Z_113) );
  XNOR2_X1 U2326 ( .A(key_in[113]), .B(data_in[113]), .ZN(n5122) );
  OAI22_X1 U2327 ( .A1(n5414), .A2(n4477), .B1(n5123), .B2(n5409), .ZN(
        U49_Z_112) );
  XNOR2_X1 U2328 ( .A(key_in[112]), .B(data_in[112]), .ZN(n5123) );
  OAI22_X1 U2329 ( .A1(n5416), .A2(n4478), .B1(n5124), .B2(n5409), .ZN(
        U49_Z_111) );
  XNOR2_X1 U2330 ( .A(key_in[111]), .B(data_in[111]), .ZN(n5124) );
  OAI22_X1 U2331 ( .A1(n5419), .A2(n4479), .B1(n5125), .B2(n5409), .ZN(
        U49_Z_110) );
  XNOR2_X1 U2332 ( .A(key_in[110]), .B(data_in[110]), .ZN(n5125) );
  OAI22_X1 U2333 ( .A1(n5415), .A2(n4480), .B1(n5127), .B2(n5409), .ZN(
        U49_Z_109) );
  XNOR2_X1 U2334 ( .A(key_in[109]), .B(data_in[109]), .ZN(n5127) );
  OAI22_X1 U2335 ( .A1(n5419), .A2(n4481), .B1(n5128), .B2(n5409), .ZN(
        U49_Z_108) );
  XNOR2_X1 U2336 ( .A(key_in[108]), .B(data_in[108]), .ZN(n5128) );
  OAI22_X1 U2337 ( .A1(n5417), .A2(n4482), .B1(n5129), .B2(n5409), .ZN(
        U49_Z_107) );
  XNOR2_X1 U2338 ( .A(key_in[107]), .B(data_in[107]), .ZN(n5129) );
  OAI22_X1 U2339 ( .A1(n5419), .A2(n4483), .B1(n5130), .B2(n5409), .ZN(
        U49_Z_106) );
  XNOR2_X1 U2340 ( .A(key_in[106]), .B(data_in[106]), .ZN(n5130) );
  OAI22_X1 U2341 ( .A1(n5415), .A2(n4484), .B1(n5131), .B2(n5410), .ZN(
        U49_Z_105) );
  XNOR2_X1 U2342 ( .A(key_in[105]), .B(data_in[105]), .ZN(n5131) );
  OAI22_X1 U2343 ( .A1(n5418), .A2(n4485), .B1(n5132), .B2(n5412), .ZN(
        U49_Z_104) );
  XNOR2_X1 U2344 ( .A(key_in[104]), .B(data_in[104]), .ZN(n5132) );
  OAI22_X1 U2345 ( .A1(n5417), .A2(n4486), .B1(n5133), .B2(n5413), .ZN(
        U49_Z_103) );
  XNOR2_X1 U2346 ( .A(key_in[103]), .B(data_in[103]), .ZN(n5133) );
  OAI22_X1 U2347 ( .A1(n5419), .A2(n4487), .B1(n5134), .B2(n5411), .ZN(
        U49_Z_102) );
  XNOR2_X1 U2348 ( .A(key_in[102]), .B(data_in[102]), .ZN(n5134) );
  OAI22_X1 U2349 ( .A1(n5419), .A2(n4488), .B1(n5135), .B2(n5409), .ZN(
        U49_Z_101) );
  XNOR2_X1 U2350 ( .A(key_in[101]), .B(data_in[101]), .ZN(n5135) );
  OAI22_X1 U2351 ( .A1(n5414), .A2(n4489), .B1(n5136), .B2(n5012), .ZN(
        U49_Z_100) );
  XNOR2_X1 U2352 ( .A(key_in[100]), .B(data_in[100]), .ZN(n5136) );
  OAI22_X1 U2353 ( .A1(n5414), .A2(n4577), .B1(n5115), .B2(n5410), .ZN(
        U49_Z_12) );
  XNOR2_X1 U2354 ( .A(key_in[12]), .B(data_in[12]), .ZN(n5115) );
  OAI22_X1 U2355 ( .A1(n5419), .A2(n4578), .B1(n5126), .B2(n5409), .ZN(
        U49_Z_11) );
  XNOR2_X1 U2356 ( .A(key_in[11]), .B(data_in[11]), .ZN(n5126) );
  OAI22_X1 U2357 ( .A1(n5417), .A2(n4579), .B1(n5137), .B2(n5410), .ZN(
        U49_Z_10) );
  XNOR2_X1 U2358 ( .A(key_in[10]), .B(data_in[10]), .ZN(n5137) );
  OAI22_X1 U2359 ( .A1(n5417), .A2(n4588), .B1(n5138), .B2(n5412), .ZN(U49_Z_1) );
  XNOR2_X1 U2360 ( .A(key_in[1]), .B(data_in[1]), .ZN(n5138) );
  OAI22_X1 U2361 ( .A1(n5418), .A2(n4589), .B1(n5139), .B2(n5413), .ZN(U49_Z_0) );
  XNOR2_X1 U2362 ( .A(key_in[0]), .B(data_in[0]), .ZN(n5139) );
  OAI22_X1 U2363 ( .A1(n5415), .A2(n4517), .B1(n5041), .B2(n5413), .ZN(
        U49_Z_72) );
  XNOR2_X1 U2364 ( .A(key_in[72]), .B(data_in[72]), .ZN(n5041) );
  OAI22_X1 U2365 ( .A1(n5414), .A2(n4518), .B1(n5042), .B2(n5410), .ZN(
        U49_Z_71) );
  XNOR2_X1 U2366 ( .A(key_in[71]), .B(data_in[71]), .ZN(n5042) );
  OAI22_X1 U2367 ( .A1(n5417), .A2(n4519), .B1(n5043), .B2(n5409), .ZN(
        U49_Z_70) );
  XNOR2_X1 U2368 ( .A(key_in[70]), .B(data_in[70]), .ZN(n5043) );
  OAI22_X1 U2369 ( .A1(n5415), .A2(n4520), .B1(n5045), .B2(n5411), .ZN(
        U49_Z_69) );
  XNOR2_X1 U2370 ( .A(key_in[69]), .B(data_in[69]), .ZN(n5045) );
  OAI22_X1 U2371 ( .A1(n5419), .A2(n4521), .B1(n5046), .B2(n5412), .ZN(
        U49_Z_68) );
  XNOR2_X1 U2372 ( .A(key_in[68]), .B(data_in[68]), .ZN(n5046) );
  OAI22_X1 U2373 ( .A1(n5418), .A2(n4522), .B1(n5047), .B2(n5413), .ZN(
        U49_Z_67) );
  XNOR2_X1 U2374 ( .A(key_in[67]), .B(data_in[67]), .ZN(n5047) );
  OAI22_X1 U2375 ( .A1(n5417), .A2(n4523), .B1(n5048), .B2(n5411), .ZN(
        U49_Z_66) );
  XNOR2_X1 U2376 ( .A(key_in[66]), .B(data_in[66]), .ZN(n5048) );
  OAI22_X1 U2377 ( .A1(n5417), .A2(n4524), .B1(n5049), .B2(n5412), .ZN(
        U49_Z_65) );
  XNOR2_X1 U2378 ( .A(key_in[65]), .B(data_in[65]), .ZN(n5049) );
  OAI22_X1 U2379 ( .A1(n5416), .A2(n4525), .B1(n5050), .B2(n5411), .ZN(
        U49_Z_64) );
  XNOR2_X1 U2380 ( .A(key_in[64]), .B(data_in[64]), .ZN(n5050) );
  OAI22_X1 U2381 ( .A1(n5414), .A2(n4526), .B1(n5051), .B2(n5413), .ZN(
        U49_Z_63) );
  XNOR2_X1 U2382 ( .A(key_in[63]), .B(data_in[63]), .ZN(n5051) );
  OAI22_X1 U2383 ( .A1(n5416), .A2(n4527), .B1(n5052), .B2(n5409), .ZN(
        U49_Z_62) );
  XNOR2_X1 U2384 ( .A(key_in[62]), .B(data_in[62]), .ZN(n5052) );
  OAI22_X1 U2385 ( .A1(n5419), .A2(n4528), .B1(n5053), .B2(n5410), .ZN(
        U49_Z_61) );
  XNOR2_X1 U2386 ( .A(key_in[61]), .B(data_in[61]), .ZN(n5053) );
  OAI22_X1 U2387 ( .A1(n5417), .A2(n4529), .B1(n5054), .B2(n5409), .ZN(
        U49_Z_60) );
  XNOR2_X1 U2388 ( .A(key_in[60]), .B(data_in[60]), .ZN(n5054) );
  OAI22_X1 U2389 ( .A1(n5415), .A2(n4530), .B1(n5056), .B2(n5409), .ZN(
        U49_Z_59) );
  XNOR2_X1 U2390 ( .A(key_in[59]), .B(data_in[59]), .ZN(n5056) );
  OAI22_X1 U2391 ( .A1(n5414), .A2(n4531), .B1(n5057), .B2(n5012), .ZN(
        U49_Z_58) );
  XNOR2_X1 U2392 ( .A(key_in[58]), .B(data_in[58]), .ZN(n5057) );
  OAI22_X1 U2393 ( .A1(n5415), .A2(n4532), .B1(n5058), .B2(n5412), .ZN(
        U49_Z_57) );
  XNOR2_X1 U2394 ( .A(key_in[57]), .B(data_in[57]), .ZN(n5058) );
  OAI22_X1 U2395 ( .A1(n5417), .A2(n4533), .B1(n5059), .B2(n5409), .ZN(
        U49_Z_56) );
  XNOR2_X1 U2396 ( .A(key_in[56]), .B(data_in[56]), .ZN(n5059) );
  OAI22_X1 U2397 ( .A1(n5416), .A2(n4534), .B1(n5060), .B2(n5410), .ZN(
        U49_Z_55) );
  XNOR2_X1 U2398 ( .A(key_in[55]), .B(data_in[55]), .ZN(n5060) );
  OAI22_X1 U2399 ( .A1(n5414), .A2(n4535), .B1(n5061), .B2(n5412), .ZN(
        U49_Z_54) );
  XNOR2_X1 U2400 ( .A(key_in[54]), .B(data_in[54]), .ZN(n5061) );
  OAI22_X1 U2401 ( .A1(n5418), .A2(n4536), .B1(n5062), .B2(n5413), .ZN(
        U49_Z_53) );
  XNOR2_X1 U2402 ( .A(key_in[53]), .B(data_in[53]), .ZN(n5062) );
  OAI22_X1 U2403 ( .A1(n5417), .A2(n4537), .B1(n5063), .B2(n5411), .ZN(
        U49_Z_52) );
  XNOR2_X1 U2404 ( .A(key_in[52]), .B(data_in[52]), .ZN(n5063) );
  OAI22_X1 U2405 ( .A1(n5418), .A2(n4538), .B1(n5064), .B2(n5411), .ZN(
        U49_Z_51) );
  XNOR2_X1 U2406 ( .A(key_in[51]), .B(data_in[51]), .ZN(n5064) );
  OAI22_X1 U2407 ( .A1(n5418), .A2(n4539), .B1(n5065), .B2(n5411), .ZN(
        U49_Z_50) );
  XNOR2_X1 U2408 ( .A(key_in[50]), .B(data_in[50]), .ZN(n5065) );
  OAI22_X1 U2409 ( .A1(n5415), .A2(n4540), .B1(n5067), .B2(n5410), .ZN(
        U49_Z_49) );
  XNOR2_X1 U2410 ( .A(key_in[49]), .B(data_in[49]), .ZN(n5067) );
  OAI22_X1 U2411 ( .A1(n5417), .A2(n4541), .B1(n5068), .B2(n5411), .ZN(
        U49_Z_48) );
  XNOR2_X1 U2412 ( .A(key_in[48]), .B(data_in[48]), .ZN(n5068) );
  OAI22_X1 U2413 ( .A1(n5418), .A2(n4542), .B1(n5069), .B2(n5410), .ZN(
        U49_Z_47) );
  XNOR2_X1 U2414 ( .A(key_in[47]), .B(data_in[47]), .ZN(n5069) );
  OAI22_X1 U2415 ( .A1(n5414), .A2(n4543), .B1(n5070), .B2(n5409), .ZN(
        U49_Z_46) );
  XNOR2_X1 U2416 ( .A(key_in[46]), .B(data_in[46]), .ZN(n5070) );
  OAI22_X1 U2417 ( .A1(n5415), .A2(n4544), .B1(n5071), .B2(n5412), .ZN(
        U49_Z_45) );
  XNOR2_X1 U2418 ( .A(key_in[45]), .B(data_in[45]), .ZN(n5071) );
  OAI22_X1 U2419 ( .A1(n5414), .A2(n4545), .B1(n5072), .B2(n5412), .ZN(
        U49_Z_44) );
  XNOR2_X1 U2420 ( .A(key_in[44]), .B(data_in[44]), .ZN(n5072) );
  OAI22_X1 U2421 ( .A1(n5418), .A2(n4546), .B1(n5073), .B2(n5413), .ZN(
        U49_Z_43) );
  XNOR2_X1 U2422 ( .A(key_in[43]), .B(data_in[43]), .ZN(n5073) );
  OAI22_X1 U2423 ( .A1(n5414), .A2(n4547), .B1(n5074), .B2(n5411), .ZN(
        U49_Z_42) );
  XNOR2_X1 U2424 ( .A(key_in[42]), .B(data_in[42]), .ZN(n5074) );
  OAI22_X1 U2425 ( .A1(n5415), .A2(n4548), .B1(n5075), .B2(n5410), .ZN(
        U49_Z_41) );
  XNOR2_X1 U2426 ( .A(key_in[41]), .B(data_in[41]), .ZN(n5075) );
  OAI22_X1 U2427 ( .A1(n5418), .A2(n4549), .B1(n5076), .B2(n5409), .ZN(
        U49_Z_40) );
  XNOR2_X1 U2428 ( .A(key_in[40]), .B(data_in[40]), .ZN(n5076) );
  OAI22_X1 U2429 ( .A1(n5417), .A2(n4550), .B1(n5078), .B2(n5012), .ZN(
        U49_Z_39) );
  XNOR2_X1 U2430 ( .A(key_in[39]), .B(data_in[39]), .ZN(n5078) );
  OAI22_X1 U2431 ( .A1(n5419), .A2(n4551), .B1(n5079), .B2(n5012), .ZN(
        U49_Z_38) );
  XNOR2_X1 U2432 ( .A(key_in[38]), .B(data_in[38]), .ZN(n5079) );
  OAI22_X1 U2433 ( .A1(n5415), .A2(n4552), .B1(n5080), .B2(n5012), .ZN(
        U49_Z_37) );
  XNOR2_X1 U2434 ( .A(key_in[37]), .B(data_in[37]), .ZN(n5080) );
  OAI22_X1 U2435 ( .A1(n5418), .A2(n4553), .B1(n5081), .B2(n5012), .ZN(
        U49_Z_36) );
  XNOR2_X1 U2436 ( .A(key_in[36]), .B(data_in[36]), .ZN(n5081) );
  OAI22_X1 U2437 ( .A1(n5415), .A2(n4554), .B1(n5082), .B2(n5012), .ZN(
        U49_Z_35) );
  XNOR2_X1 U2438 ( .A(key_in[35]), .B(data_in[35]), .ZN(n5082) );
  OAI22_X1 U2439 ( .A1(n5414), .A2(n4555), .B1(n5083), .B2(n5012), .ZN(
        U49_Z_34) );
  XNOR2_X1 U2440 ( .A(key_in[34]), .B(data_in[34]), .ZN(n5083) );
  OAI22_X1 U2441 ( .A1(n5415), .A2(n4556), .B1(n5084), .B2(n5410), .ZN(
        U49_Z_33) );
  XNOR2_X1 U2442 ( .A(key_in[33]), .B(data_in[33]), .ZN(n5084) );
  OAI22_X1 U2443 ( .A1(n5417), .A2(n4557), .B1(n5085), .B2(n5409), .ZN(
        U49_Z_32) );
  XNOR2_X1 U2444 ( .A(key_in[32]), .B(data_in[32]), .ZN(n5085) );
  OAI22_X1 U2445 ( .A1(n5417), .A2(n4558), .B1(n5086), .B2(n5012), .ZN(
        U49_Z_31) );
  XNOR2_X1 U2446 ( .A(key_in[31]), .B(data_in[31]), .ZN(n5086) );
  OAI22_X1 U2447 ( .A1(n5417), .A2(n4559), .B1(n5087), .B2(n5012), .ZN(
        U49_Z_30) );
  XNOR2_X1 U2448 ( .A(key_in[30]), .B(data_in[30]), .ZN(n5087) );
  OAI22_X1 U2449 ( .A1(n5417), .A2(n4560), .B1(n5089), .B2(n5012), .ZN(
        U49_Z_29) );
  XNOR2_X1 U2450 ( .A(key_in[29]), .B(data_in[29]), .ZN(n5089) );
  OAI22_X1 U2451 ( .A1(n5418), .A2(n4561), .B1(n5090), .B2(n5012), .ZN(
        U49_Z_28) );
  XNOR2_X1 U2452 ( .A(key_in[28]), .B(data_in[28]), .ZN(n5090) );
  OAI22_X1 U2453 ( .A1(n5416), .A2(n4562), .B1(n5091), .B2(n5012), .ZN(
        U49_Z_27) );
  XNOR2_X1 U2454 ( .A(key_in[27]), .B(data_in[27]), .ZN(n5091) );
  OAI22_X1 U2455 ( .A1(n5419), .A2(n4563), .B1(n5092), .B2(n5012), .ZN(
        U49_Z_26) );
  XNOR2_X1 U2456 ( .A(key_in[26]), .B(data_in[26]), .ZN(n5092) );
  OAI22_X1 U2457 ( .A1(n5416), .A2(n4564), .B1(n5093), .B2(n5012), .ZN(
        U49_Z_25) );
  XNOR2_X1 U2458 ( .A(key_in[25]), .B(data_in[25]), .ZN(n5093) );
  OAI22_X1 U2459 ( .A1(n5419), .A2(n4565), .B1(n5094), .B2(n5012), .ZN(
        U49_Z_24) );
  XNOR2_X1 U2460 ( .A(key_in[24]), .B(data_in[24]), .ZN(n5094) );
  OAI22_X1 U2461 ( .A1(n5418), .A2(n4582), .B1(n5044), .B2(n5410), .ZN(U49_Z_7) );
  XNOR2_X1 U2462 ( .A(key_in[7]), .B(data_in[7]), .ZN(n5044) );
  OAI22_X1 U2463 ( .A1(n5419), .A2(n4583), .B1(n5055), .B2(n5413), .ZN(U49_Z_6) );
  XNOR2_X1 U2464 ( .A(key_in[6]), .B(data_in[6]), .ZN(n5055) );
  OAI22_X1 U2465 ( .A1(n5419), .A2(n4584), .B1(n5066), .B2(n5410), .ZN(U49_Z_5) );
  XNOR2_X1 U2466 ( .A(key_in[5]), .B(data_in[5]), .ZN(n5066) );
  OAI22_X1 U2467 ( .A1(n5414), .A2(n4585), .B1(n5077), .B2(n5012), .ZN(U49_Z_4) );
  XNOR2_X1 U2468 ( .A(key_in[4]), .B(data_in[4]), .ZN(n5077) );
  OAI22_X1 U2469 ( .A1(n5417), .A2(n4586), .B1(n5088), .B2(n5012), .ZN(U49_Z_3) );
  XNOR2_X1 U2470 ( .A(key_in[3]), .B(data_in[3]), .ZN(n5088) );
  NAND2_X1 U2471 ( .A1(n4595), .A2(r424_A_0_), .ZN(n5009) );
  OR3_X1 U2472 ( .A1(n4597), .A2(n3261), .A3(n4592), .ZN(n5141) );
  INV_X1 U2473 ( .A(n5145), .ZN(n4591) );
  OAI21_X1 U2474 ( .B1(n4598), .B2(n4874), .A(n4873), .ZN(n5145) );
  INV_X1 U2475 ( .A(n4878), .ZN(n4358) );
  AOI22_X1 U2476 ( .A1(n5423), .A2(U99_DATA1_99), .B1(n5427), .B2(key_in[99]), 
        .ZN(n4878) );
  INV_X1 U2477 ( .A(n4880), .ZN(n4359) );
  AOI22_X1 U2478 ( .A1(n5423), .A2(U99_DATA1_98), .B1(n5429), .B2(key_in[98]), 
        .ZN(n4880) );
  INV_X1 U2479 ( .A(n4881), .ZN(n4360) );
  AOI22_X1 U2480 ( .A1(n5420), .A2(U99_DATA1_97), .B1(n5430), .B2(key_in[97]), 
        .ZN(n4881) );
  INV_X1 U2481 ( .A(n4882), .ZN(n4361) );
  AOI22_X1 U2482 ( .A1(n4879), .A2(U99_DATA1_96), .B1(n5426), .B2(key_in[96]), 
        .ZN(n4882) );
  INV_X1 U2483 ( .A(n4883), .ZN(n4362) );
  AOI22_X1 U2484 ( .A1(n5424), .A2(U99_DATA1_95), .B1(n5429), .B2(key_in[95]), 
        .ZN(n4883) );
  INV_X1 U2485 ( .A(n4884), .ZN(n4363) );
  AOI22_X1 U2486 ( .A1(n5422), .A2(U99_DATA1_94), .B1(n5429), .B2(key_in[94]), 
        .ZN(n4884) );
  INV_X1 U2487 ( .A(n4885), .ZN(n4364) );
  AOI22_X1 U2488 ( .A1(n5421), .A2(U99_DATA1_93), .B1(n5426), .B2(key_in[93]), 
        .ZN(n4885) );
  INV_X1 U2489 ( .A(n4886), .ZN(n4365) );
  AOI22_X1 U2490 ( .A1(n5423), .A2(U99_DATA1_92), .B1(n5430), .B2(key_in[92]), 
        .ZN(n4886) );
  INV_X1 U2491 ( .A(n4975), .ZN(n4331) );
  AOI22_X1 U2492 ( .A1(n5423), .A2(U99_DATA1_126), .B1(n5427), .B2(key_in[126]), .ZN(n4975) );
  INV_X1 U2493 ( .A(n4976), .ZN(n4332) );
  AOI22_X1 U2494 ( .A1(n5423), .A2(U99_DATA1_125), .B1(n5425), .B2(key_in[125]), .ZN(n4976) );
  INV_X1 U2495 ( .A(n4977), .ZN(n4333) );
  AOI22_X1 U2496 ( .A1(n5423), .A2(U99_DATA1_124), .B1(n5430), .B2(key_in[124]), .ZN(n4977) );
  INV_X1 U2497 ( .A(n4978), .ZN(n4334) );
  AOI22_X1 U2498 ( .A1(n5423), .A2(U99_DATA1_123), .B1(n5425), .B2(key_in[123]), .ZN(n4978) );
  INV_X1 U2499 ( .A(n4979), .ZN(n4335) );
  AOI22_X1 U2500 ( .A1(n5423), .A2(U99_DATA1_122), .B1(n5428), .B2(key_in[122]), .ZN(n4979) );
  INV_X1 U2501 ( .A(n4980), .ZN(n4336) );
  AOI22_X1 U2502 ( .A1(n5423), .A2(U99_DATA1_121), .B1(n5426), .B2(key_in[121]), .ZN(n4980) );
  INV_X1 U2503 ( .A(n4981), .ZN(n4337) );
  AOI22_X1 U2504 ( .A1(n5423), .A2(U99_DATA1_120), .B1(n5425), .B2(key_in[120]), .ZN(n4981) );
  INV_X1 U2505 ( .A(n4983), .ZN(n4338) );
  AOI22_X1 U2506 ( .A1(n5422), .A2(U99_DATA1_119), .B1(n5427), .B2(key_in[119]), .ZN(n4983) );
  INV_X1 U2507 ( .A(n4984), .ZN(n4339) );
  AOI22_X1 U2508 ( .A1(n5422), .A2(U99_DATA1_118), .B1(n5427), .B2(key_in[118]), .ZN(n4984) );
  INV_X1 U2509 ( .A(n4985), .ZN(n4340) );
  AOI22_X1 U2510 ( .A1(n5422), .A2(U99_DATA1_117), .B1(n5427), .B2(key_in[117]), .ZN(n4985) );
  INV_X1 U2511 ( .A(n4986), .ZN(n4341) );
  AOI22_X1 U2512 ( .A1(n5422), .A2(U99_DATA1_116), .B1(n5427), .B2(key_in[116]), .ZN(n4986) );
  INV_X1 U2513 ( .A(n4987), .ZN(n4342) );
  AOI22_X1 U2514 ( .A1(n5422), .A2(U99_DATA1_115), .B1(n5426), .B2(key_in[115]), .ZN(n4987) );
  INV_X1 U2515 ( .A(n4988), .ZN(n4343) );
  AOI22_X1 U2516 ( .A1(n5422), .A2(U99_DATA1_114), .B1(n5426), .B2(key_in[114]), .ZN(n4988) );
  INV_X1 U2517 ( .A(n4989), .ZN(n4344) );
  AOI22_X1 U2518 ( .A1(n5422), .A2(U99_DATA1_113), .B1(n5426), .B2(key_in[113]), .ZN(n4989) );
  INV_X1 U2519 ( .A(n4990), .ZN(n4345) );
  AOI22_X1 U2520 ( .A1(n5422), .A2(U99_DATA1_112), .B1(n5426), .B2(key_in[112]), .ZN(n4990) );
  INV_X1 U2521 ( .A(n4991), .ZN(n4346) );
  AOI22_X1 U2522 ( .A1(n5422), .A2(U99_DATA1_111), .B1(n5426), .B2(key_in[111]), .ZN(n4991) );
  INV_X1 U2523 ( .A(n4992), .ZN(n4347) );
  AOI22_X1 U2524 ( .A1(n5422), .A2(U99_DATA1_110), .B1(n5425), .B2(key_in[110]), .ZN(n4992) );
  INV_X1 U2525 ( .A(n4994), .ZN(n4348) );
  AOI22_X1 U2526 ( .A1(n5422), .A2(U99_DATA1_109), .B1(n5425), .B2(key_in[109]), .ZN(n4994) );
  INV_X1 U2527 ( .A(n4995), .ZN(n4349) );
  AOI22_X1 U2528 ( .A1(n5421), .A2(U99_DATA1_108), .B1(n5425), .B2(key_in[108]), .ZN(n4995) );
  INV_X1 U2529 ( .A(n4996), .ZN(n4350) );
  AOI22_X1 U2530 ( .A1(n5421), .A2(U99_DATA1_107), .B1(n5425), .B2(key_in[107]), .ZN(n4996) );
  INV_X1 U2531 ( .A(n4997), .ZN(n4351) );
  AOI22_X1 U2532 ( .A1(n5421), .A2(U99_DATA1_106), .B1(n5429), .B2(key_in[106]), .ZN(n4997) );
  INV_X1 U2533 ( .A(n4998), .ZN(n4352) );
  AOI22_X1 U2534 ( .A1(n5421), .A2(U99_DATA1_105), .B1(n5425), .B2(key_in[105]), .ZN(n4998) );
  INV_X1 U2535 ( .A(n4999), .ZN(n4353) );
  AOI22_X1 U2536 ( .A1(n5421), .A2(U99_DATA1_104), .B1(n5428), .B2(key_in[104]), .ZN(n4999) );
  INV_X1 U2537 ( .A(n5000), .ZN(n4354) );
  AOI22_X1 U2538 ( .A1(n5421), .A2(U99_DATA1_103), .B1(n5427), .B2(key_in[103]), .ZN(n5000) );
  INV_X1 U2539 ( .A(n5001), .ZN(n4355) );
  AOI22_X1 U2540 ( .A1(n5421), .A2(U99_DATA1_102), .B1(n5426), .B2(key_in[102]), .ZN(n5001) );
  INV_X1 U2541 ( .A(n5002), .ZN(n4356) );
  AOI22_X1 U2542 ( .A1(n5421), .A2(U99_DATA1_101), .B1(n5428), .B2(key_in[101]), .ZN(n5002) );
  INV_X1 U2543 ( .A(n5003), .ZN(n4357) );
  AOI22_X1 U2544 ( .A1(n5421), .A2(U99_DATA1_100), .B1(n5426), .B2(key_in[100]), .ZN(n5003) );
  INV_X1 U2545 ( .A(n4887), .ZN(n4366) );
  AOI22_X1 U2546 ( .A1(n5421), .A2(U99_DATA1_91), .B1(n5425), .B2(key_in[91]), 
        .ZN(n4887) );
  INV_X1 U2547 ( .A(n4888), .ZN(n4367) );
  AOI22_X1 U2548 ( .A1(n5424), .A2(U99_DATA1_90), .B1(n5430), .B2(key_in[90]), 
        .ZN(n4888) );
  INV_X1 U2549 ( .A(n4890), .ZN(n4368) );
  AOI22_X1 U2550 ( .A1(n5421), .A2(U99_DATA1_89), .B1(n5427), .B2(key_in[89]), 
        .ZN(n4890) );
  INV_X1 U2551 ( .A(n4891), .ZN(n4369) );
  AOI22_X1 U2552 ( .A1(n5422), .A2(U99_DATA1_88), .B1(n5425), .B2(key_in[88]), 
        .ZN(n4891) );
  INV_X1 U2553 ( .A(n4892), .ZN(n4370) );
  AOI22_X1 U2554 ( .A1(n5421), .A2(U99_DATA1_87), .B1(n5425), .B2(key_in[87]), 
        .ZN(n4892) );
  INV_X1 U2555 ( .A(n4893), .ZN(n4371) );
  AOI22_X1 U2556 ( .A1(n5423), .A2(U99_DATA1_86), .B1(n5426), .B2(key_in[86]), 
        .ZN(n4893) );
  INV_X1 U2557 ( .A(n4894), .ZN(n4372) );
  AOI22_X1 U2558 ( .A1(n5420), .A2(U99_DATA1_85), .B1(n5429), .B2(key_in[85]), 
        .ZN(n4894) );
  INV_X1 U2559 ( .A(n4895), .ZN(n4373) );
  AOI22_X1 U2560 ( .A1(n4879), .A2(U99_DATA1_84), .B1(n5426), .B2(key_in[84]), 
        .ZN(n4895) );
  INV_X1 U2561 ( .A(n4896), .ZN(n4374) );
  AOI22_X1 U2562 ( .A1(n5424), .A2(U99_DATA1_83), .B1(n5429), .B2(key_in[83]), 
        .ZN(n4896) );
  INV_X1 U2563 ( .A(n4897), .ZN(n4375) );
  AOI22_X1 U2564 ( .A1(n5422), .A2(U99_DATA1_82), .B1(n5430), .B2(key_in[82]), 
        .ZN(n4897) );
  INV_X1 U2565 ( .A(n4898), .ZN(n4376) );
  AOI22_X1 U2566 ( .A1(n4879), .A2(U99_DATA1_81), .B1(n5429), .B2(key_in[81]), 
        .ZN(n4898) );
  INV_X1 U2567 ( .A(n4899), .ZN(n4377) );
  AOI22_X1 U2568 ( .A1(n5423), .A2(U99_DATA1_80), .B1(n5428), .B2(key_in[80]), 
        .ZN(n4899) );
  INV_X1 U2569 ( .A(n4901), .ZN(n4378) );
  AOI22_X1 U2570 ( .A1(n5422), .A2(U99_DATA1_79), .B1(n5427), .B2(key_in[79]), 
        .ZN(n4901) );
  INV_X1 U2571 ( .A(n4902), .ZN(n4379) );
  AOI22_X1 U2572 ( .A1(n5420), .A2(U99_DATA1_78), .B1(n5425), .B2(key_in[78]), 
        .ZN(n4902) );
  INV_X1 U2573 ( .A(n4903), .ZN(n4380) );
  AOI22_X1 U2574 ( .A1(n4879), .A2(U99_DATA1_77), .B1(n5430), .B2(key_in[77]), 
        .ZN(n4903) );
  INV_X1 U2575 ( .A(n4904), .ZN(n4381) );
  AOI22_X1 U2576 ( .A1(n5420), .A2(U99_DATA1_76), .B1(n5430), .B2(key_in[76]), 
        .ZN(n4904) );
  INV_X1 U2577 ( .A(n4905), .ZN(n4382) );
  AOI22_X1 U2578 ( .A1(n5424), .A2(U99_DATA1_75), .B1(n5428), .B2(key_in[75]), 
        .ZN(n4905) );
  INV_X1 U2579 ( .A(n4906), .ZN(n4383) );
  AOI22_X1 U2580 ( .A1(n5424), .A2(U99_DATA1_74), .B1(n5429), .B2(key_in[74]), 
        .ZN(n4906) );
  INV_X1 U2581 ( .A(n4907), .ZN(n4384) );
  AOI22_X1 U2582 ( .A1(n5422), .A2(U99_DATA1_73), .B1(n5426), .B2(key_in[73]), 
        .ZN(n4907) );
  INV_X1 U2583 ( .A(n4908), .ZN(n4385) );
  AOI22_X1 U2584 ( .A1(n5421), .A2(U99_DATA1_72), .B1(n5427), .B2(key_in[72]), 
        .ZN(n4908) );
  INV_X1 U2585 ( .A(n4909), .ZN(n4386) );
  AOI22_X1 U2586 ( .A1(n5423), .A2(U99_DATA1_71), .B1(n5425), .B2(key_in[71]), 
        .ZN(n4909) );
  INV_X1 U2587 ( .A(n4910), .ZN(n4387) );
  AOI22_X1 U2588 ( .A1(n5420), .A2(U99_DATA1_70), .B1(n5426), .B2(key_in[70]), 
        .ZN(n4910) );
  INV_X1 U2589 ( .A(n4912), .ZN(n4388) );
  AOI22_X1 U2590 ( .A1(n5420), .A2(U99_DATA1_69), .B1(n5428), .B2(key_in[69]), 
        .ZN(n4912) );
  INV_X1 U2591 ( .A(n4913), .ZN(n4389) );
  AOI22_X1 U2592 ( .A1(n4879), .A2(U99_DATA1_68), .B1(n5427), .B2(key_in[68]), 
        .ZN(n4913) );
  INV_X1 U2593 ( .A(n4914), .ZN(n4390) );
  AOI22_X1 U2594 ( .A1(n4879), .A2(U99_DATA1_67), .B1(n5427), .B2(key_in[67]), 
        .ZN(n4914) );
  INV_X1 U2595 ( .A(n4915), .ZN(n4391) );
  AOI22_X1 U2596 ( .A1(n5420), .A2(U99_DATA1_66), .B1(n5430), .B2(key_in[66]), 
        .ZN(n4915) );
  INV_X1 U2597 ( .A(n4916), .ZN(n4392) );
  AOI22_X1 U2598 ( .A1(n4879), .A2(U99_DATA1_65), .B1(n5428), .B2(key_in[65]), 
        .ZN(n4916) );
  INV_X1 U2599 ( .A(n4917), .ZN(n4393) );
  AOI22_X1 U2600 ( .A1(n5424), .A2(U99_DATA1_64), .B1(n5426), .B2(key_in[64]), 
        .ZN(n4917) );
  INV_X1 U2601 ( .A(n4918), .ZN(n4394) );
  AOI22_X1 U2602 ( .A1(n5420), .A2(U99_DATA1_63), .B1(n5430), .B2(key_in[63]), 
        .ZN(n4918) );
  INV_X1 U2603 ( .A(n4919), .ZN(n4395) );
  AOI22_X1 U2604 ( .A1(n4879), .A2(U99_DATA1_62), .B1(n5428), .B2(key_in[62]), 
        .ZN(n4919) );
  INV_X1 U2605 ( .A(n4920), .ZN(n4396) );
  AOI22_X1 U2606 ( .A1(n5422), .A2(U99_DATA1_61), .B1(n5430), .B2(key_in[61]), 
        .ZN(n4920) );
  INV_X1 U2607 ( .A(n4921), .ZN(n4397) );
  AOI22_X1 U2608 ( .A1(n5420), .A2(U99_DATA1_60), .B1(n5430), .B2(key_in[60]), 
        .ZN(n4921) );
  INV_X1 U2609 ( .A(n4923), .ZN(n4398) );
  AOI22_X1 U2610 ( .A1(n5420), .A2(U99_DATA1_59), .B1(n5429), .B2(key_in[59]), 
        .ZN(n4923) );
  INV_X1 U2611 ( .A(n4924), .ZN(n4399) );
  AOI22_X1 U2612 ( .A1(n4879), .A2(U99_DATA1_58), .B1(n5429), .B2(key_in[58]), 
        .ZN(n4924) );
  INV_X1 U2613 ( .A(n4925), .ZN(n4400) );
  AOI22_X1 U2614 ( .A1(n5420), .A2(U99_DATA1_57), .B1(n5429), .B2(key_in[57]), 
        .ZN(n4925) );
  INV_X1 U2615 ( .A(n4926), .ZN(n4401) );
  AOI22_X1 U2616 ( .A1(n4879), .A2(U99_DATA1_56), .B1(n5429), .B2(key_in[56]), 
        .ZN(n4926) );
  INV_X1 U2617 ( .A(n4927), .ZN(n4402) );
  AOI22_X1 U2618 ( .A1(n5420), .A2(U99_DATA1_55), .B1(n5429), .B2(key_in[55]), 
        .ZN(n4927) );
  INV_X1 U2619 ( .A(n4928), .ZN(n4403) );
  AOI22_X1 U2620 ( .A1(n4879), .A2(U99_DATA1_54), .B1(n5428), .B2(key_in[54]), 
        .ZN(n4928) );
  INV_X1 U2621 ( .A(n4929), .ZN(n4404) );
  AOI22_X1 U2622 ( .A1(n5420), .A2(U99_DATA1_53), .B1(n5425), .B2(key_in[53]), 
        .ZN(n4929) );
  INV_X1 U2623 ( .A(n4930), .ZN(n4405) );
  AOI22_X1 U2624 ( .A1(n4879), .A2(U99_DATA1_52), .B1(n5426), .B2(key_in[52]), 
        .ZN(n4930) );
  INV_X1 U2625 ( .A(n4931), .ZN(n4406) );
  AOI22_X1 U2626 ( .A1(n5420), .A2(U99_DATA1_51), .B1(n5426), .B2(key_in[51]), 
        .ZN(n4931) );
  INV_X1 U2627 ( .A(n4932), .ZN(n4407) );
  AOI22_X1 U2628 ( .A1(n4879), .A2(U99_DATA1_50), .B1(n5428), .B2(key_in[50]), 
        .ZN(n4932) );
  INV_X1 U2629 ( .A(n4934), .ZN(n4408) );
  AOI22_X1 U2630 ( .A1(n5420), .A2(U99_DATA1_49), .B1(n5427), .B2(key_in[49]), 
        .ZN(n4934) );
  INV_X1 U2631 ( .A(n4935), .ZN(n4409) );
  AOI22_X1 U2632 ( .A1(n5424), .A2(U99_DATA1_48), .B1(n5425), .B2(key_in[48]), 
        .ZN(n4935) );
  INV_X1 U2633 ( .A(n4936), .ZN(n4410) );
  AOI22_X1 U2634 ( .A1(n5424), .A2(U99_DATA1_47), .B1(n5430), .B2(key_in[47]), 
        .ZN(n4936) );
  INV_X1 U2635 ( .A(n4937), .ZN(n4411) );
  AOI22_X1 U2636 ( .A1(n5424), .A2(U99_DATA1_46), .B1(n5428), .B2(key_in[46]), 
        .ZN(n4937) );
  INV_X1 U2637 ( .A(n4938), .ZN(n4412) );
  AOI22_X1 U2638 ( .A1(n5424), .A2(U99_DATA1_45), .B1(n5428), .B2(key_in[45]), 
        .ZN(n4938) );
  INV_X1 U2639 ( .A(n4939), .ZN(n4413) );
  AOI22_X1 U2640 ( .A1(n5424), .A2(U99_DATA1_44), .B1(n5428), .B2(key_in[44]), 
        .ZN(n4939) );
  INV_X1 U2641 ( .A(n4940), .ZN(n4414) );
  AOI22_X1 U2642 ( .A1(n5424), .A2(U99_DATA1_43), .B1(n5428), .B2(key_in[43]), 
        .ZN(n4940) );
  INV_X1 U2643 ( .A(n4941), .ZN(n4415) );
  AOI22_X1 U2644 ( .A1(n5424), .A2(U99_DATA1_42), .B1(n5428), .B2(key_in[42]), 
        .ZN(n4941) );
  INV_X1 U2645 ( .A(n4942), .ZN(n4416) );
  AOI22_X1 U2646 ( .A1(n5424), .A2(U99_DATA1_41), .B1(n5429), .B2(key_in[41]), 
        .ZN(n4942) );
  INV_X1 U2647 ( .A(n4943), .ZN(n4417) );
  AOI22_X1 U2648 ( .A1(n5424), .A2(U99_DATA1_40), .B1(n5430), .B2(key_in[40]), 
        .ZN(n4943) );
  INV_X1 U2649 ( .A(n4945), .ZN(n4418) );
  AOI22_X1 U2650 ( .A1(n5424), .A2(U99_DATA1_39), .B1(n5426), .B2(key_in[39]), 
        .ZN(n4945) );
  INV_X1 U2651 ( .A(n4946), .ZN(n4419) );
  AOI22_X1 U2652 ( .A1(n5424), .A2(U99_DATA1_38), .B1(n5429), .B2(key_in[38]), 
        .ZN(n4946) );
  INV_X1 U2653 ( .A(n4947), .ZN(n4420) );
  AOI22_X1 U2654 ( .A1(n5420), .A2(U99_DATA1_37), .B1(n5427), .B2(key_in[37]), 
        .ZN(n4947) );
  INV_X1 U2655 ( .A(n4948), .ZN(n4421) );
  AOI22_X1 U2656 ( .A1(n4879), .A2(U99_DATA1_36), .B1(n5429), .B2(key_in[36]), 
        .ZN(n4948) );
  INV_X1 U2657 ( .A(n4949), .ZN(n4422) );
  AOI22_X1 U2658 ( .A1(n5424), .A2(U99_DATA1_35), .B1(n5428), .B2(key_in[35]), 
        .ZN(n4949) );
  INV_X1 U2659 ( .A(n4950), .ZN(n4423) );
  AOI22_X1 U2660 ( .A1(n5422), .A2(U99_DATA1_34), .B1(n5427), .B2(key_in[34]), 
        .ZN(n4950) );
  INV_X1 U2661 ( .A(n4951), .ZN(n4424) );
  AOI22_X1 U2662 ( .A1(n5421), .A2(U99_DATA1_33), .B1(n5429), .B2(key_in[33]), 
        .ZN(n4951) );
  INV_X1 U2663 ( .A(n4952), .ZN(n4425) );
  AOI22_X1 U2664 ( .A1(n5423), .A2(U99_DATA1_32), .B1(n5425), .B2(key_in[32]), 
        .ZN(n4952) );
  INV_X1 U2665 ( .A(n4953), .ZN(n4426) );
  AOI22_X1 U2666 ( .A1(n5420), .A2(U99_DATA1_31), .B1(n5428), .B2(key_in[31]), 
        .ZN(n4953) );
  INV_X1 U2667 ( .A(n4954), .ZN(n4427) );
  AOI22_X1 U2668 ( .A1(n5421), .A2(U99_DATA1_30), .B1(n5430), .B2(key_in[30]), 
        .ZN(n4954) );
  INV_X1 U2669 ( .A(n4956), .ZN(n4428) );
  AOI22_X1 U2670 ( .A1(n5420), .A2(U99_DATA1_29), .B1(n5427), .B2(key_in[29]), 
        .ZN(n4956) );
  INV_X1 U2671 ( .A(n4957), .ZN(n4429) );
  AOI22_X1 U2672 ( .A1(n4879), .A2(U99_DATA1_28), .B1(n5426), .B2(key_in[28]), 
        .ZN(n4957) );
  INV_X1 U2673 ( .A(n4958), .ZN(n4430) );
  AOI22_X1 U2674 ( .A1(n5424), .A2(U99_DATA1_27), .B1(n5426), .B2(key_in[27]), 
        .ZN(n4958) );
  INV_X1 U2675 ( .A(n4959), .ZN(n4431) );
  AOI22_X1 U2676 ( .A1(n5421), .A2(U99_DATA1_26), .B1(n5427), .B2(key_in[26]), 
        .ZN(n4959) );
  INV_X1 U2677 ( .A(n4960), .ZN(n4432) );
  AOI22_X1 U2678 ( .A1(n5423), .A2(U99_DATA1_25), .B1(n5428), .B2(key_in[25]), 
        .ZN(n4960) );
  INV_X1 U2679 ( .A(n4961), .ZN(n4433) );
  AOI22_X1 U2680 ( .A1(n5420), .A2(U99_DATA1_24), .B1(n5430), .B2(key_in[24]), 
        .ZN(n4961) );
  INV_X1 U2681 ( .A(n4962), .ZN(n4434) );
  AOI22_X1 U2682 ( .A1(n4879), .A2(U99_DATA1_23), .B1(n5428), .B2(key_in[23]), 
        .ZN(n4962) );
  INV_X1 U2683 ( .A(n4963), .ZN(n4435) );
  AOI22_X1 U2684 ( .A1(n5424), .A2(U99_DATA1_22), .B1(n5425), .B2(key_in[22]), 
        .ZN(n4963) );
  INV_X1 U2685 ( .A(n4964), .ZN(n4436) );
  AOI22_X1 U2686 ( .A1(n5422), .A2(U99_DATA1_21), .B1(n5426), .B2(key_in[21]), 
        .ZN(n4964) );
  INV_X1 U2687 ( .A(n4965), .ZN(n4437) );
  AOI22_X1 U2688 ( .A1(n5421), .A2(U99_DATA1_20), .B1(n5429), .B2(key_in[20]), 
        .ZN(n4965) );
  INV_X1 U2689 ( .A(n4967), .ZN(n4438) );
  AOI22_X1 U2690 ( .A1(n5423), .A2(U99_DATA1_19), .B1(n5429), .B2(key_in[19]), 
        .ZN(n4967) );
  INV_X1 U2691 ( .A(n4968), .ZN(n4439) );
  AOI22_X1 U2692 ( .A1(n5420), .A2(U99_DATA1_18), .B1(n5426), .B2(key_in[18]), 
        .ZN(n4968) );
  INV_X1 U2693 ( .A(n4969), .ZN(n4440) );
  AOI22_X1 U2694 ( .A1(n4879), .A2(U99_DATA1_17), .B1(n5429), .B2(key_in[17]), 
        .ZN(n4969) );
  INV_X1 U2695 ( .A(n4970), .ZN(n4441) );
  AOI22_X1 U2696 ( .A1(n5424), .A2(U99_DATA1_16), .B1(n5427), .B2(key_in[16]), 
        .ZN(n4970) );
  INV_X1 U2697 ( .A(n4971), .ZN(n4442) );
  AOI22_X1 U2698 ( .A1(n5423), .A2(U99_DATA1_15), .B1(n5425), .B2(key_in[15]), 
        .ZN(n4971) );
  INV_X1 U2699 ( .A(n4972), .ZN(n4443) );
  AOI22_X1 U2700 ( .A1(n5423), .A2(U99_DATA1_14), .B1(n5430), .B2(key_in[14]), 
        .ZN(n4972) );
  INV_X1 U2701 ( .A(n4973), .ZN(n4444) );
  AOI22_X1 U2702 ( .A1(n5423), .A2(U99_DATA1_13), .B1(n5425), .B2(key_in[13]), 
        .ZN(n4973) );
  INV_X1 U2703 ( .A(n4982), .ZN(n4445) );
  AOI22_X1 U2704 ( .A1(n5423), .A2(U99_DATA1_12), .B1(n5427), .B2(key_in[12]), 
        .ZN(n4982) );
  INV_X1 U2705 ( .A(n4993), .ZN(n4446) );
  AOI22_X1 U2706 ( .A1(n5422), .A2(U99_DATA1_11), .B1(n5425), .B2(key_in[11]), 
        .ZN(n4993) );
  INV_X1 U2707 ( .A(n5004), .ZN(n4447) );
  AOI22_X1 U2708 ( .A1(n5421), .A2(U99_DATA1_10), .B1(n5429), .B2(key_in[10]), 
        .ZN(n5004) );
  INV_X1 U2709 ( .A(n4889), .ZN(n4448) );
  AOI22_X1 U2710 ( .A1(n5423), .A2(U99_DATA1_9), .B1(n5430), .B2(key_in[9]), 
        .ZN(n4889) );
  INV_X1 U2711 ( .A(n4900), .ZN(n4449) );
  AOI22_X1 U2712 ( .A1(n4879), .A2(U99_DATA1_8), .B1(n5428), .B2(key_in[8]), 
        .ZN(n4900) );
  INV_X1 U2713 ( .A(n4911), .ZN(n4450) );
  AOI22_X1 U2714 ( .A1(n4879), .A2(U99_DATA1_7), .B1(n5429), .B2(key_in[7]), 
        .ZN(n4911) );
  INV_X1 U2715 ( .A(n4922), .ZN(n4451) );
  AOI22_X1 U2716 ( .A1(n5421), .A2(U99_DATA1_6), .B1(n5429), .B2(key_in[6]), 
        .ZN(n4922) );
  INV_X1 U2717 ( .A(n4933), .ZN(n4452) );
  AOI22_X1 U2718 ( .A1(n4879), .A2(U99_DATA1_5), .B1(n5428), .B2(key_in[5]), 
        .ZN(n4933) );
  INV_X1 U2719 ( .A(n4944), .ZN(n4453) );
  AOI22_X1 U2720 ( .A1(n5424), .A2(U99_DATA1_4), .B1(n5428), .B2(key_in[4]), 
        .ZN(n4944) );
  INV_X1 U2721 ( .A(n4955), .ZN(n4454) );
  AOI22_X1 U2722 ( .A1(n5422), .A2(U99_DATA1_3), .B1(n5426), .B2(key_in[3]), 
        .ZN(n4955) );
  INV_X1 U2723 ( .A(n4966), .ZN(n4455) );
  AOI22_X1 U2724 ( .A1(n5422), .A2(U99_DATA1_2), .B1(n5427), .B2(key_in[2]), 
        .ZN(n4966) );
  INV_X1 U2725 ( .A(n5005), .ZN(n4456) );
  AOI22_X1 U2726 ( .A1(n5421), .A2(U99_DATA1_1), .B1(n5427), .B2(key_in[1]), 
        .ZN(n5005) );
  INV_X1 U2727 ( .A(n5006), .ZN(n4457) );
  AOI22_X1 U2728 ( .A1(n5421), .A2(U99_DATA1_0), .B1(n5425), .B2(key_in[0]), 
        .ZN(n5006) );
  INV_X1 U2729 ( .A(n4974), .ZN(n4330) );
  AOI22_X1 U2730 ( .A1(n5423), .A2(U99_DATA1_127), .B1(n5428), .B2(key_in[127]), .ZN(n4974) );
  INV_X1 U2731 ( .A(n5463), .ZN(n5457) );
  CLKBUF_X1 U2732 ( .A(n5471), .Z(n5465) );
  CLKBUF_X1 U2733 ( .A(n5464), .Z(n5466) );
  CLKBUF_X1 U2734 ( .A(n5464), .Z(n5467) );
  CLKBUF_X1 U2735 ( .A(n5464), .Z(n5468) );
  CLKBUF_X1 U2736 ( .A(n5464), .Z(n5469) );
  CLKBUF_X1 U2737 ( .A(n5464), .Z(n5470) );
  CLKBUF_X1 U2738 ( .A(n5464), .Z(n5471) );
  CLKBUF_X1 U2739 ( .A(U47_Z_1), .Z(n5472) );
  CLKBUF_X1 U2740 ( .A(U47_Z_1), .Z(n5473) );
  CLKBUF_X1 U2741 ( .A(n5472), .Z(n5474) );
  CLKBUF_X1 U2742 ( .A(n5472), .Z(n5475) );
  AOI21_X2 U1348 ( .B1(n4593), .B2(n5143), .A(ready), .ZN(U46_Z_1) );
  NAND3_X2 U1349 ( .A1(n3262), .A2(n5408), .A3(n4730), .ZN(n4602) );
  OAI21_X2 U1350 ( .B1(n4868), .B2(n4201), .A(n4730), .ZN(n4733) );
  CLKBUF_X2 U1352 ( .A(n5444), .Z(n5449) );
  CLKBUF_X2 U1353 ( .A(n5445), .Z(n5448) );
  CLKBUF_X2 U1360 ( .A(n5417), .Z(n5415) );
  CLKBUF_X2 U1362 ( .A(n5463), .Z(n5458) );
  CLKBUF_X2 U1381 ( .A(n5463), .Z(n5459) );
  CLKBUF_X2 U1384 ( .A(n5463), .Z(n5461) );
  CLKBUF_X2 U1385 ( .A(n5463), .Z(n5460) );
  CLKBUF_X2 U1386 ( .A(n5418), .Z(n5417) );
  CLKBUF_X2 U1387 ( .A(n5419), .Z(n5418) );
  INV_X2 U1397 ( .A(n5012), .ZN(n5419) );
  CLKBUF_X2 U1398 ( .A(n5447), .Z(n5451) );
  CLKBUF_X2 U1399 ( .A(n4601), .Z(n5454) );
  NAND2_X2 U1404 ( .A1(n4730), .A2(n4201), .ZN(n4601) );
  CLKBUF_X2 U1409 ( .A(n5431), .Z(n5441) );
  CLKBUF_X2 U1580 ( .A(n4733), .Z(n5431) );
  CLKBUF_X1 U2213 ( .A(n4602), .Z(n5443) );
  CLKBUF_X2 U2743 ( .A(n4602), .Z(n5447) );
  CLKBUF_X2 R2_U1123 ( .A(R2_n2343), .Z(R2_n2353) );
  CLKBUF_X2 R2_U1122 ( .A(R2_n1811), .Z(R2_n2376) );
  CLKBUF_X2 R2_U1120 ( .A(R2_n2376), .Z(R2_n2375) );
  CLKBUF_X2 R2_U1119 ( .A(R2_n2398), .Z(R2_n2401) );
  CLKBUF_X2 R2_U1118 ( .A(R2_n2398), .Z(R2_n2402) );
  CLKBUF_X2 R2_U1117 ( .A(R2_n2398), .Z(R2_n2404) );
  CLKBUF_X2 R2_U1116 ( .A(R2_n2398), .Z(R2_n2403) );
  AND2_X2 R2_U1113 ( .A1(R2_n2336), .A2(R2_n1807), .ZN(R2_U23_Z_1) );
  CLKBUF_X2 R2_U1108 ( .A(R2_U23_Z_1), .Z(R2_n2398) );
  NAND2_X2 R2_U1107 ( .A1(R2_n2333), .A2(R2_n2334), .ZN(R2_n2071) );
  CLKBUF_X2 R2_U1106 ( .A(R2_n2071), .Z(R2_n2361) );
  CLKBUF_X2 R2_U1105 ( .A(R2_n1802), .Z(R2_n2386) );
  CLKBUF_X2 R2_U1061 ( .A(R2_n2386), .Z(R2_n2387) );
  CLKBUF_X2 R2_U332 ( .A(R2_n2386), .Z(R2_n2388) );
  CLKBUF_X2 R2_U64 ( .A(R2_n2386), .Z(R2_n2389) );
  CLKBUF_X2 R2_U61 ( .A(R2_n2386), .Z(R2_n2390) );
  NAND4_X2 R2_U60 ( .A1(R2_n1515), .A2(R2_n2337), .A3(R2_n2334), .A4(R2_n1805), 
        .ZN(R2_n2200) );
  CLKBUF_X2 R2_U54 ( .A(R2_n2200), .Z(R2_n2343) );
  CLKBUF_X2 R2_U53 ( .A(R2_n1940), .Z(R2_n2373) );
  CLKBUF_X2 R2_U52 ( .A(R2_n2371), .Z(R2_n2374) );
  NAND2_X2 R2_U49 ( .A1(R2_n2334), .A2(R2_n2336), .ZN(R2_n1811) );
  AND2_X2 R2_U42 ( .A1(R2_n2069), .A2(R2_n610), .ZN(R2_n1941) );
  CLKBUF_X2 R2_U24 ( .A(R2_n1941), .Z(R2_n2365) );
  CLKBUF_X2 R2_U23 ( .A(R2_U22_Z_1), .Z(R2_n2395) );
  CLKBUF_X2 R2_U20 ( .A(R2_n2395), .Z(R2_n2396) );
  CLKBUF_X2 R2_U18 ( .A(R2_n2403), .Z(R2_n2400) );
  CLKBUF_X2 R2_U17 ( .A(R2_U24_Z_1), .Z(R2_n2406) );
  CLKBUF_X2 R2_U14 ( .A(R2_n2406), .Z(R2_n2407) );
  AND3_X2 R2_U12 ( .A1(R2_n1805), .A2(R2_n1807), .A3(R2_n2337), .ZN(R2_U24_Z_1) );
  NOR2_X2 R2_U8 ( .A1(R2_n1802), .A2(R2_n610), .ZN(R2_n1940) );
  AND2_X2 R2_U7 ( .A1(R2_n2333), .A2(R2_n1807), .ZN(R2_U22_Z_1) );
  NOR3_X2 R2_U6 ( .A1(n3391), .A2(n3262), .A3(R2_n2335), .ZN(R2_U21_Z_1) );
  CLKBUF_X1 R2_U1121 ( .A(R2_U24_Z_1), .Z(R2_n2405) );
  CLKBUF_X1 R2_U1115 ( .A(R2_n2403), .Z(R2_n2399) );
  CLKBUF_X1 R2_U1114 ( .A(R2_n2395), .Z(R2_n2397) );
  CLKBUF_X1 R2_U1112 ( .A(R2_n2391), .Z(R2_n2394) );
  CLKBUF_X1 R2_U1111 ( .A(R2_U21_Z_1), .Z(R2_n2393) );
  CLKBUF_X1 R2_U1110 ( .A(R2_n2393), .Z(R2_n2392) );
  CLKBUF_X1 R2_U1109 ( .A(R2_U21_Z_1), .Z(R2_n2391) );
  AOI22_X1 R2_U1104 ( .A1(R2_n2355), .A2(R2_n1281), .B1(R2_n2362), .B2(
        R2_U16_DATA1_23), .ZN(R2_n2175) );
  INV_X1 R2_U1103 ( .A(R2_n2175), .ZN(R2_n154) );
  AOI22_X1 R2_U1102 ( .A1(R2_n2360), .A2(R2_n1282), .B1(R2_n2363), .B2(
        R2_U16_DATA1_24), .ZN(R2_n2174) );
  INV_X1 R2_U1101 ( .A(R2_n2174), .ZN(R2_n155) );
  AOI22_X1 R2_U1100 ( .A1(R2_n2357), .A2(R2_n1283), .B1(R2_n2364), .B2(
        R2_U16_DATA1_25), .ZN(R2_n2173) );
  INV_X1 R2_U1099 ( .A(R2_n2173), .ZN(R2_n156) );
  AOI22_X1 R2_U1098 ( .A1(R2_n2357), .A2(R2_n1284), .B1(R2_n2362), .B2(
        R2_U16_DATA1_26), .ZN(R2_n2172) );
  INV_X1 R2_U1097 ( .A(R2_n2172), .ZN(R2_n157) );
  AOI22_X1 R2_U1096 ( .A1(R2_n2359), .A2(R2_n1285), .B1(R2_n2364), .B2(
        R2_U16_DATA1_27), .ZN(R2_n2171) );
  INV_X1 R2_U1095 ( .A(R2_n2171), .ZN(R2_n158) );
  AOI22_X1 R2_U1094 ( .A1(R2_n2358), .A2(R2_n1286), .B1(R2_n2363), .B2(
        R2_U16_DATA1_28), .ZN(R2_n2170) );
  INV_X1 R2_U1093 ( .A(R2_n2170), .ZN(R2_n159) );
  AOI22_X1 R2_U1092 ( .A1(R2_n2357), .A2(R2_n1287), .B1(R2_n2364), .B2(
        R2_U16_DATA1_29), .ZN(R2_n2169) );
  INV_X1 R2_U1091 ( .A(R2_n2169), .ZN(R2_n160) );
  AOI22_X1 R2_U1090 ( .A1(R2_n2357), .A2(R2_n1288), .B1(R2_n2362), .B2(
        R2_U16_DATA1_30), .ZN(R2_n2168) );
  INV_X1 R2_U1089 ( .A(R2_n2168), .ZN(R2_n161) );
  AOI22_X1 R2_U1088 ( .A1(R2_n2356), .A2(R2_n1289), .B1(R2_n2363), .B2(
        R2_U16_DATA1_31), .ZN(R2_n2167) );
  INV_X1 R2_U1087 ( .A(R2_n2167), .ZN(R2_n162) );
  AOI22_X1 R2_U1086 ( .A1(R2_n2355), .A2(R2_n1290), .B1(R2_n2364), .B2(
        R2_U16_DATA1_32), .ZN(R2_n2166) );
  INV_X1 R2_U1085 ( .A(R2_n2166), .ZN(R2_n163) );
  AOI22_X1 R2_U1084 ( .A1(R2_n2356), .A2(R2_n1291), .B1(R2_n2361), .B2(
        R2_U16_DATA1_33), .ZN(R2_n2165) );
  INV_X1 R2_U1083 ( .A(R2_n2165), .ZN(R2_n164) );
  AOI22_X1 R2_U1082 ( .A1(R2_n2356), .A2(R2_n1292), .B1(R2_n2361), .B2(
        R2_U16_DATA1_34), .ZN(R2_n2164) );
  INV_X1 R2_U1081 ( .A(R2_n2164), .ZN(R2_n165) );
  AOI22_X1 R2_U1080 ( .A1(R2_n2360), .A2(R2_n1293), .B1(R2_n2361), .B2(
        R2_U16_DATA1_35), .ZN(R2_n2163) );
  INV_X1 R2_U1079 ( .A(R2_n2163), .ZN(R2_n166) );
  AOI22_X1 R2_U1078 ( .A1(R2_n2360), .A2(R2_n1294), .B1(R2_n2361), .B2(
        R2_U16_DATA1_36), .ZN(R2_n2162) );
  INV_X1 R2_U1077 ( .A(R2_n2162), .ZN(R2_n167) );
  AOI22_X1 R2_U1076 ( .A1(R2_n2359), .A2(R2_n1295), .B1(R2_n2361), .B2(
        R2_U16_DATA1_37), .ZN(R2_n2161) );
  INV_X1 R2_U1075 ( .A(R2_n2161), .ZN(R2_n168) );
  AOI22_X1 R2_U1074 ( .A1(R2_n2358), .A2(R2_n1296), .B1(R2_n2364), .B2(
        R2_U16_DATA1_38), .ZN(R2_n2160) );
  INV_X1 R2_U1073 ( .A(R2_n2160), .ZN(R2_n169) );
  AOI22_X1 R2_U1072 ( .A1(R2_n2357), .A2(R2_n1297), .B1(R2_n2362), .B2(
        R2_U16_DATA1_39), .ZN(R2_n2159) );
  INV_X1 R2_U1071 ( .A(R2_n2159), .ZN(R2_n170) );
  AOI22_X1 R2_U1070 ( .A1(R2_n2355), .A2(R2_n1298), .B1(R2_n2364), .B2(
        R2_U16_DATA1_40), .ZN(R2_n2158) );
  INV_X1 R2_U1069 ( .A(R2_n2158), .ZN(R2_n171) );
  AOI22_X1 R2_U1068 ( .A1(R2_n2356), .A2(R2_n1299), .B1(R2_n2362), .B2(
        R2_U16_DATA1_41), .ZN(R2_n2157) );
  INV_X1 R2_U1067 ( .A(R2_n2157), .ZN(R2_n172) );
  AOI22_X1 R2_U1066 ( .A1(R2_n2359), .A2(R2_n1300), .B1(R2_n2363), .B2(
        R2_U16_DATA1_42), .ZN(R2_n2156) );
  INV_X1 R2_U1065 ( .A(R2_n2156), .ZN(R2_n173) );
  AOI22_X1 R2_U1064 ( .A1(R2_n2359), .A2(R2_n1301), .B1(R2_n2364), .B2(
        R2_U16_DATA1_43), .ZN(R2_n2155) );
  INV_X1 R2_U1063 ( .A(R2_n2155), .ZN(R2_n174) );
  AOI22_X1 R2_U1062 ( .A1(R2_n2358), .A2(R2_n1302), .B1(R2_n2364), .B2(
        R2_U16_DATA1_44), .ZN(R2_n2154) );
  INV_X1 R2_U1057 ( .A(R2_n2154), .ZN(R2_n175) );
  AOI22_X1 R2_U1056 ( .A1(R2_n2357), .A2(R2_n1303), .B1(R2_n2362), .B2(
        R2_U16_DATA1_45), .ZN(R2_n2153) );
  INV_X1 R2_U1055 ( .A(R2_n2153), .ZN(R2_n176) );
  AOI22_X1 R2_U1054 ( .A1(R2_n2356), .A2(R2_n1304), .B1(R2_n2362), .B2(
        R2_U16_DATA1_46), .ZN(R2_n2152) );
  INV_X1 R2_U1053 ( .A(R2_n2152), .ZN(R2_n177) );
  AOI22_X1 R2_U1052 ( .A1(R2_n2355), .A2(R2_n1305), .B1(R2_n2363), .B2(
        R2_U16_DATA1_47), .ZN(R2_n2151) );
  INV_X1 R2_U1051 ( .A(R2_n2151), .ZN(R2_n178) );
  AOI22_X1 R2_U1050 ( .A1(R2_n2360), .A2(R2_n1306), .B1(R2_n2364), .B2(
        R2_U16_DATA1_48), .ZN(R2_n2150) );
  INV_X1 R2_U1049 ( .A(R2_n2150), .ZN(R2_n179) );
  AOI22_X1 R2_U1048 ( .A1(R2_n2359), .A2(R2_n1307), .B1(R2_n2361), .B2(
        R2_U16_DATA1_49), .ZN(R2_n2149) );
  INV_X1 R2_U1047 ( .A(R2_n2149), .ZN(R2_n180) );
  AOI22_X1 R2_U1046 ( .A1(R2_n2358), .A2(R2_n1308), .B1(R2_n2362), .B2(
        R2_U16_DATA1_50), .ZN(R2_n2148) );
  INV_X1 R2_U1045 ( .A(R2_n2148), .ZN(R2_n181) );
  AOI22_X1 R2_U1044 ( .A1(R2_n2357), .A2(R2_n1309), .B1(R2_n2361), .B2(
        R2_U16_DATA1_51), .ZN(R2_n2147) );
  INV_X1 R2_U1043 ( .A(R2_n2147), .ZN(R2_n182) );
  AOI22_X1 R2_U1042 ( .A1(R2_n2356), .A2(R2_n1310), .B1(R2_n2362), .B2(
        R2_U16_DATA1_52), .ZN(R2_n2146) );
  INV_X1 R2_U1041 ( .A(R2_n2146), .ZN(R2_n183) );
  AOI22_X1 R2_U1040 ( .A1(R2_n2355), .A2(R2_n1311), .B1(R2_n2361), .B2(
        R2_U16_DATA1_53), .ZN(R2_n2145) );
  INV_X1 R2_U1039 ( .A(R2_n2145), .ZN(R2_n184) );
  AOI22_X1 R2_U1038 ( .A1(R2_n2360), .A2(R2_n1312), .B1(R2_n2363), .B2(
        R2_U16_DATA1_54), .ZN(R2_n2144) );
  INV_X1 R2_U1037 ( .A(R2_n2144), .ZN(R2_n185) );
  AOI22_X1 R2_U1036 ( .A1(R2_n2359), .A2(R2_n1313), .B1(R2_n2361), .B2(
        R2_U16_DATA1_55), .ZN(R2_n2143) );
  INV_X1 R2_U1035 ( .A(R2_n2143), .ZN(R2_n186) );
  AOI22_X1 R2_U1034 ( .A1(R2_n2359), .A2(R2_n1314), .B1(R2_n2362), .B2(
        R2_U16_DATA1_56), .ZN(R2_n2142) );
  INV_X1 R2_U1033 ( .A(R2_n2142), .ZN(R2_n187) );
  AOI22_X1 R2_U1032 ( .A1(R2_n2359), .A2(R2_n1315), .B1(R2_n2364), .B2(
        R2_U16_DATA1_57), .ZN(R2_n2141) );
  INV_X1 R2_U1031 ( .A(R2_n2141), .ZN(R2_n188) );
  AOI22_X1 R2_U1030 ( .A1(R2_n2359), .A2(R2_n1316), .B1(R2_n2354), .B2(
        R2_U16_DATA1_58), .ZN(R2_n2140) );
  INV_X1 R2_U1029 ( .A(R2_n2140), .ZN(R2_n189) );
  AOI22_X1 R2_U1028 ( .A1(R2_n2359), .A2(R2_n1317), .B1(R2_n2354), .B2(
        R2_U16_DATA1_59), .ZN(R2_n2139) );
  INV_X1 R2_U1027 ( .A(R2_n2139), .ZN(R2_n190) );
  AOI22_X1 R2_U1026 ( .A1(R2_n2359), .A2(R2_n1318), .B1(R2_n2364), .B2(
        R2_U16_DATA1_60), .ZN(R2_n2138) );
  INV_X1 R2_U1025 ( .A(R2_n2138), .ZN(R2_n191) );
  AOI22_X1 R2_U1024 ( .A1(R2_n2359), .A2(R2_n1319), .B1(R2_n2361), .B2(
        R2_U16_DATA1_61), .ZN(R2_n2137) );
  INV_X1 R2_U1023 ( .A(R2_n2137), .ZN(R2_n192) );
  AOI22_X1 R2_U1022 ( .A1(R2_n2359), .A2(R2_n1320), .B1(R2_n2071), .B2(
        R2_U16_DATA1_62), .ZN(R2_n2136) );
  INV_X1 R2_U1021 ( .A(R2_n2136), .ZN(R2_n193) );
  AOI22_X1 R2_U1020 ( .A1(R2_n2359), .A2(R2_n1321), .B1(R2_n2362), .B2(
        R2_U16_DATA1_63), .ZN(R2_n2135) );
  INV_X1 R2_U1019 ( .A(R2_n2135), .ZN(R2_n194) );
  AOI22_X1 R2_U1018 ( .A1(R2_n2359), .A2(R2_n1322), .B1(R2_n2354), .B2(
        R2_U16_DATA1_64), .ZN(R2_n2134) );
  INV_X1 R2_U1017 ( .A(R2_n2134), .ZN(R2_n195) );
  AOI22_X1 R2_U1016 ( .A1(R2_n2359), .A2(R2_n1323), .B1(R2_n2361), .B2(
        R2_U16_DATA1_65), .ZN(R2_n2133) );
  INV_X1 R2_U1015 ( .A(R2_n2133), .ZN(R2_n196) );
  AOI22_X1 R2_U1014 ( .A1(R2_n2359), .A2(R2_n1324), .B1(R2_n2361), .B2(
        R2_U16_DATA1_66), .ZN(R2_n2132) );
  INV_X1 R2_U1013 ( .A(R2_n2132), .ZN(R2_n197) );
  AOI22_X1 R2_U1012 ( .A1(R2_n2359), .A2(R2_n1325), .B1(R2_n2363), .B2(
        R2_U16_DATA1_67), .ZN(R2_n2131) );
  INV_X1 R2_U1011 ( .A(R2_n2131), .ZN(R2_n198) );
  AOI22_X1 R2_U1010 ( .A1(R2_n2358), .A2(R2_n1326), .B1(R2_n2361), .B2(
        R2_U16_DATA1_68), .ZN(R2_n2130) );
  INV_X1 R2_U1009 ( .A(R2_n2130), .ZN(R2_n199) );
  AOI22_X1 R2_U1008 ( .A1(R2_n2358), .A2(R2_n1327), .B1(R2_n2362), .B2(
        R2_U16_DATA1_69), .ZN(R2_n2129) );
  INV_X1 R2_U1007 ( .A(R2_n2129), .ZN(R2_n200) );
  AOI22_X1 R2_U1006 ( .A1(R2_n2358), .A2(R2_n1328), .B1(R2_n2364), .B2(
        R2_U16_DATA1_70), .ZN(R2_n2128) );
  INV_X1 R2_U1005 ( .A(R2_n2128), .ZN(R2_n201) );
  AOI22_X1 R2_U1004 ( .A1(R2_n2358), .A2(R2_n1329), .B1(R2_n2361), .B2(
        R2_U16_DATA1_71), .ZN(R2_n2127) );
  INV_X1 R2_U1003 ( .A(R2_n2127), .ZN(R2_n202) );
  AOI22_X1 R2_U1002 ( .A1(R2_n2358), .A2(R2_n1330), .B1(R2_n2362), .B2(
        R2_U16_DATA1_72), .ZN(R2_n2126) );
  INV_X1 R2_U1001 ( .A(R2_n2126), .ZN(R2_n203) );
  AOI22_X1 R2_U1000 ( .A1(R2_n2358), .A2(R2_n1331), .B1(R2_n2361), .B2(
        R2_U16_DATA1_73), .ZN(R2_n2125) );
  INV_X1 R2_U999 ( .A(R2_n2125), .ZN(R2_n204) );
  AOI22_X1 R2_U998 ( .A1(R2_n2358), .A2(R2_n1332), .B1(R2_n2361), .B2(
        R2_U16_DATA1_74), .ZN(R2_n2124) );
  INV_X1 R2_U997 ( .A(R2_n2124), .ZN(R2_n205) );
  AOI22_X1 R2_U996 ( .A1(R2_n2358), .A2(R2_n1333), .B1(R2_n2071), .B2(
        R2_U16_DATA1_75), .ZN(R2_n2123) );
  INV_X1 R2_U995 ( .A(R2_n2123), .ZN(R2_n206) );
  AOI22_X1 R2_U994 ( .A1(R2_n2358), .A2(R2_n1334), .B1(R2_n2071), .B2(
        R2_U16_DATA1_76), .ZN(R2_n2122) );
  INV_X1 R2_U993 ( .A(R2_n2122), .ZN(R2_n207) );
  AOI22_X1 R2_U992 ( .A1(R2_n2358), .A2(R2_n1335), .B1(R2_n2361), .B2(
        R2_U16_DATA1_77), .ZN(R2_n2121) );
  INV_X1 R2_U991 ( .A(R2_n2121), .ZN(R2_n208) );
  AOI22_X1 R2_U990 ( .A1(R2_n2358), .A2(R2_n1336), .B1(R2_n2071), .B2(
        R2_U16_DATA1_78), .ZN(R2_n2120) );
  INV_X1 R2_U989 ( .A(R2_n2120), .ZN(R2_n209) );
  AOI22_X1 R2_U988 ( .A1(R2_n2358), .A2(R2_n1337), .B1(R2_n2363), .B2(
        R2_U16_DATA1_79), .ZN(R2_n2119) );
  INV_X1 R2_U987 ( .A(R2_n2119), .ZN(R2_n210) );
  AOI22_X1 R2_U986 ( .A1(R2_n2357), .A2(R2_n1338), .B1(R2_n2361), .B2(
        R2_U16_DATA1_80), .ZN(R2_n2118) );
  INV_X1 R2_U985 ( .A(R2_n2118), .ZN(R2_n211) );
  AOI22_X1 R2_U984 ( .A1(R2_n2357), .A2(R2_n1339), .B1(R2_n2361), .B2(
        R2_U16_DATA1_81), .ZN(R2_n2117) );
  INV_X1 R2_U983 ( .A(R2_n2117), .ZN(R2_n212) );
  AOI22_X1 R2_U982 ( .A1(R2_n2357), .A2(R2_n1340), .B1(R2_n2361), .B2(
        R2_U16_DATA1_82), .ZN(R2_n2116) );
  INV_X1 R2_U981 ( .A(R2_n2116), .ZN(R2_n213) );
  AOI22_X1 R2_U980 ( .A1(R2_n2357), .A2(R2_n1341), .B1(R2_n2361), .B2(
        R2_U16_DATA1_83), .ZN(R2_n2115) );
  INV_X1 R2_U979 ( .A(R2_n2115), .ZN(R2_n214) );
  AOI22_X1 R2_U978 ( .A1(R2_n2357), .A2(R2_n1342), .B1(R2_n2071), .B2(
        R2_U16_DATA1_84), .ZN(R2_n2114) );
  INV_X1 R2_U977 ( .A(R2_n2114), .ZN(R2_n215) );
  AOI22_X1 R2_U976 ( .A1(R2_n2357), .A2(R2_n1343), .B1(R2_n2363), .B2(
        R2_U16_DATA1_85), .ZN(R2_n2113) );
  INV_X1 R2_U975 ( .A(R2_n2113), .ZN(R2_n216) );
  AOI22_X1 R2_U974 ( .A1(R2_n2357), .A2(R2_n1344), .B1(R2_n2361), .B2(
        R2_U16_DATA1_86), .ZN(R2_n2112) );
  INV_X1 R2_U973 ( .A(R2_n2112), .ZN(R2_n217) );
  AOI22_X1 R2_U972 ( .A1(R2_n2357), .A2(R2_n1345), .B1(R2_n2364), .B2(
        R2_U16_DATA1_87), .ZN(R2_n2111) );
  INV_X1 R2_U971 ( .A(R2_n2111), .ZN(R2_n218) );
  AOI22_X1 R2_U970 ( .A1(R2_n2357), .A2(R2_n1346), .B1(R2_n2361), .B2(
        R2_U16_DATA1_88), .ZN(R2_n2110) );
  INV_X1 R2_U969 ( .A(R2_n2110), .ZN(R2_n219) );
  AOI22_X1 R2_U968 ( .A1(R2_n2357), .A2(R2_n1347), .B1(R2_n2361), .B2(
        R2_U16_DATA1_89), .ZN(R2_n2109) );
  INV_X1 R2_U967 ( .A(R2_n2109), .ZN(R2_n220) );
  AOI22_X1 R2_U966 ( .A1(R2_n2357), .A2(R2_n1348), .B1(R2_n2071), .B2(
        R2_U16_DATA1_90), .ZN(R2_n2108) );
  INV_X1 R2_U965 ( .A(R2_n2108), .ZN(R2_n221) );
  AOI22_X1 R2_U964 ( .A1(R2_n2357), .A2(R2_n1349), .B1(R2_n2071), .B2(
        R2_U16_DATA1_91), .ZN(R2_n2107) );
  INV_X1 R2_U963 ( .A(R2_n2107), .ZN(R2_n222) );
  AOI22_X1 R2_U962 ( .A1(R2_n2356), .A2(R2_n1350), .B1(R2_n2361), .B2(
        R2_U16_DATA1_92), .ZN(R2_n2106) );
  INV_X1 R2_U961 ( .A(R2_n2106), .ZN(R2_n223) );
  AOI22_X1 R2_U960 ( .A1(R2_n2355), .A2(R2_n1351), .B1(R2_n2071), .B2(
        R2_U16_DATA1_93), .ZN(R2_n2105) );
  INV_X1 R2_U959 ( .A(R2_n2105), .ZN(R2_n224) );
  AOI22_X1 R2_U958 ( .A1(R2_n2360), .A2(R2_n1352), .B1(R2_n2361), .B2(
        R2_U16_DATA1_94), .ZN(R2_n2104) );
  INV_X1 R2_U957 ( .A(R2_n2104), .ZN(R2_n353) );
  AOI22_X1 R2_U956 ( .A1(R2_n2358), .A2(R2_n1353), .B1(R2_n2361), .B2(
        R2_U16_DATA1_95), .ZN(R2_n2103) );
  INV_X1 R2_U955 ( .A(R2_n2103), .ZN(R2_n354) );
  AOI22_X1 R2_U954 ( .A1(R2_n2359), .A2(R2_n1354), .B1(R2_n2361), .B2(
        R2_U16_DATA1_96), .ZN(R2_n2102) );
  INV_X1 R2_U953 ( .A(R2_n2102), .ZN(R2_n355) );
  AOI22_X1 R2_U952 ( .A1(R2_n2358), .A2(R2_n1355), .B1(R2_n2071), .B2(
        R2_U16_DATA1_97), .ZN(R2_n2101) );
  INV_X1 R2_U951 ( .A(R2_n2101), .ZN(R2_n356) );
  AOI22_X1 R2_U950 ( .A1(R2_n2357), .A2(R2_n1356), .B1(R2_n2364), .B2(
        R2_U16_DATA1_98), .ZN(R2_n2100) );
  INV_X1 R2_U949 ( .A(R2_n2100), .ZN(R2_n357) );
  AOI22_X1 R2_U948 ( .A1(R2_n2356), .A2(R2_n1357), .B1(R2_n2362), .B2(
        R2_U16_DATA1_99), .ZN(R2_n2099) );
  INV_X1 R2_U947 ( .A(R2_n2099), .ZN(R2_n358) );
  AOI22_X1 R2_U946 ( .A1(R2_n2355), .A2(R2_n1358), .B1(R2_n2363), .B2(
        R2_U16_DATA1_100), .ZN(R2_n2098) );
  INV_X1 R2_U945 ( .A(R2_n2098), .ZN(R2_n359) );
  AOI22_X1 R2_U944 ( .A1(R2_n2360), .A2(R2_n1359), .B1(R2_n2364), .B2(
        R2_U16_DATA1_101), .ZN(R2_n2097) );
  INV_X1 R2_U943 ( .A(R2_n2097), .ZN(R2_n360) );
  AOI22_X1 R2_U942 ( .A1(R2_n2357), .A2(R2_n1360), .B1(R2_n2361), .B2(
        R2_U16_DATA1_102), .ZN(R2_n2096) );
  INV_X1 R2_U941 ( .A(R2_n2096), .ZN(R2_n361) );
  AOI22_X1 R2_U940 ( .A1(R2_n2359), .A2(R2_n1361), .B1(R2_n2363), .B2(
        R2_U16_DATA1_103), .ZN(R2_n2095) );
  INV_X1 R2_U939 ( .A(R2_n2095), .ZN(R2_n362) );
  AOI22_X1 R2_U938 ( .A1(R2_n2356), .A2(R2_n1362), .B1(R2_n2361), .B2(
        R2_U16_DATA1_104), .ZN(R2_n2094) );
  INV_X1 R2_U937 ( .A(R2_n2094), .ZN(R2_n363) );
  AOI22_X1 R2_U936 ( .A1(R2_n2356), .A2(R2_n1363), .B1(R2_n2363), .B2(
        R2_U16_DATA1_105), .ZN(R2_n2093) );
  INV_X1 R2_U935 ( .A(R2_n2093), .ZN(R2_n364) );
  AOI22_X1 R2_U934 ( .A1(R2_n2356), .A2(R2_n1364), .B1(R2_n2361), .B2(
        R2_U16_DATA1_106), .ZN(R2_n2092) );
  INV_X1 R2_U933 ( .A(R2_n2092), .ZN(R2_n365) );
  AOI22_X1 R2_U932 ( .A1(R2_n2356), .A2(R2_n1365), .B1(R2_n2361), .B2(
        R2_U16_DATA1_107), .ZN(R2_n2091) );
  INV_X1 R2_U931 ( .A(R2_n2091), .ZN(R2_n366) );
  AOI22_X1 R2_U930 ( .A1(R2_n2356), .A2(R2_n1366), .B1(R2_n2363), .B2(
        R2_U16_DATA1_108), .ZN(R2_n2090) );
  INV_X1 R2_U929 ( .A(R2_n2090), .ZN(R2_n367) );
  AOI22_X1 R2_U928 ( .A1(R2_n2356), .A2(R2_n1367), .B1(R2_n2361), .B2(
        R2_U16_DATA1_109), .ZN(R2_n2089) );
  INV_X1 R2_U927 ( .A(R2_n2089), .ZN(R2_n368) );
  AOI22_X1 R2_U926 ( .A1(R2_n2356), .A2(R2_n1368), .B1(R2_n2362), .B2(
        R2_U16_DATA1_110), .ZN(R2_n2088) );
  INV_X1 R2_U925 ( .A(R2_n2088), .ZN(R2_n369) );
  AOI22_X1 R2_U924 ( .A1(R2_n2356), .A2(R2_n1369), .B1(R2_n2361), .B2(
        R2_U16_DATA1_111), .ZN(R2_n2087) );
  INV_X1 R2_U923 ( .A(R2_n2087), .ZN(R2_n370) );
  AOI22_X1 R2_U922 ( .A1(R2_n2356), .A2(R2_n1370), .B1(R2_n2364), .B2(
        R2_U16_DATA1_112), .ZN(R2_n2086) );
  INV_X1 R2_U921 ( .A(R2_n2086), .ZN(R2_n371) );
  AOI22_X1 R2_U920 ( .A1(R2_n2356), .A2(R2_n1371), .B1(R2_n2071), .B2(
        R2_U16_DATA1_113), .ZN(R2_n2085) );
  INV_X1 R2_U919 ( .A(R2_n2085), .ZN(R2_n372) );
  AOI22_X1 R2_U918 ( .A1(R2_n2356), .A2(R2_n1372), .B1(R2_n2361), .B2(
        R2_U16_DATA1_114), .ZN(R2_n2084) );
  INV_X1 R2_U917 ( .A(R2_n2084), .ZN(R2_n373) );
  AOI22_X1 R2_U916 ( .A1(R2_n2356), .A2(R2_n1373), .B1(R2_n2071), .B2(
        R2_U16_DATA1_115), .ZN(R2_n2083) );
  INV_X1 R2_U915 ( .A(R2_n2083), .ZN(R2_n374) );
  AOI22_X1 R2_U914 ( .A1(R2_n2355), .A2(R2_n1374), .B1(R2_n2071), .B2(
        R2_U16_DATA1_116), .ZN(R2_n2082) );
  INV_X1 R2_U913 ( .A(R2_n2082), .ZN(R2_n375) );
  AOI22_X1 R2_U912 ( .A1(R2_n2355), .A2(R2_n1375), .B1(R2_n2071), .B2(
        R2_U16_DATA1_117), .ZN(R2_n2081) );
  INV_X1 R2_U911 ( .A(R2_n2081), .ZN(R2_n376) );
  AOI22_X1 R2_U910 ( .A1(R2_n2355), .A2(R2_n1376), .B1(R2_n2363), .B2(
        R2_U16_DATA1_118), .ZN(R2_n2080) );
  INV_X1 R2_U909 ( .A(R2_n2080), .ZN(R2_n377) );
  AOI22_X1 R2_U908 ( .A1(R2_n2355), .A2(R2_n1377), .B1(R2_n2361), .B2(
        R2_U16_DATA1_119), .ZN(R2_n2079) );
  INV_X1 R2_U907 ( .A(R2_n2079), .ZN(R2_n378) );
  AOI22_X1 R2_U906 ( .A1(R2_n2355), .A2(R2_n1378), .B1(R2_n2361), .B2(
        R2_U16_DATA1_120), .ZN(R2_n2078) );
  INV_X1 R2_U905 ( .A(R2_n2078), .ZN(R2_n379) );
  AOI22_X1 R2_U904 ( .A1(R2_n2355), .A2(R2_n1379), .B1(R2_n2362), .B2(
        R2_U16_DATA1_121), .ZN(R2_n2077) );
  INV_X1 R2_U903 ( .A(R2_n2077), .ZN(R2_n380) );
  AOI22_X1 R2_U902 ( .A1(R2_n2355), .A2(R2_n1380), .B1(R2_n2363), .B2(
        R2_U16_DATA1_122), .ZN(R2_n2076) );
  INV_X1 R2_U901 ( .A(R2_n2076), .ZN(R2_n381) );
  AOI22_X1 R2_U900 ( .A1(R2_n2355), .A2(R2_n1381), .B1(R2_n2361), .B2(
        R2_U16_DATA1_123), .ZN(R2_n2075) );
  INV_X1 R2_U899 ( .A(R2_n2075), .ZN(R2_n382) );
  AOI22_X1 R2_U898 ( .A1(R2_n2355), .A2(R2_n1382), .B1(R2_n2362), .B2(
        R2_U16_DATA1_124), .ZN(R2_n2074) );
  INV_X1 R2_U897 ( .A(R2_n2074), .ZN(R2_n383) );
  AOI22_X1 R2_U896 ( .A1(R2_n2355), .A2(R2_n1383), .B1(R2_n2361), .B2(
        R2_U16_DATA1_125), .ZN(R2_n2073) );
  INV_X1 R2_U895 ( .A(R2_n2073), .ZN(R2_n384) );
  AOI22_X1 R2_U894 ( .A1(R2_n2355), .A2(R2_n1384), .B1(R2_n2362), .B2(
        R2_U16_DATA1_126), .ZN(R2_n2072) );
  INV_X1 R2_U893 ( .A(R2_n2072), .ZN(R2_n385) );
  AOI22_X1 R2_U892 ( .A1(R2_n2355), .A2(R2_n1385), .B1(R2_n2364), .B2(
        R2_U16_DATA1_127), .ZN(R2_n2070) );
  INV_X1 R2_U891 ( .A(R2_n2070), .ZN(R2_n386) );
  AOI22_X1 R2_U890 ( .A1(R2_n2360), .A2(R2_n1266), .B1(R2_n2361), .B2(
        R2_U16_DATA1_8), .ZN(R2_n2190) );
  INV_X1 R2_U889 ( .A(R2_n2190), .ZN(R2_n139) );
  AOI22_X1 R2_U888 ( .A1(R2_n2360), .A2(R2_n1267), .B1(R2_n2364), .B2(
        R2_U16_DATA1_9), .ZN(R2_n2189) );
  INV_X1 R2_U887 ( .A(R2_n2189), .ZN(R2_n140) );
  AOI22_X1 R2_U886 ( .A1(R2_n2360), .A2(R2_n1268), .B1(R2_n2364), .B2(
        R2_U16_DATA1_10), .ZN(R2_n2188) );
  INV_X1 R2_U885 ( .A(R2_n2188), .ZN(R2_n141) );
  AOI22_X1 R2_U884 ( .A1(R2_n2360), .A2(R2_n1269), .B1(R2_n2364), .B2(
        R2_U16_DATA1_11), .ZN(R2_n2187) );
  INV_X1 R2_U883 ( .A(R2_n2187), .ZN(R2_n142) );
  AOI22_X1 R2_U882 ( .A1(R2_n2360), .A2(R2_n1270), .B1(R2_n2364), .B2(
        R2_U16_DATA1_12), .ZN(R2_n2186) );
  INV_X1 R2_U881 ( .A(R2_n2186), .ZN(R2_n143) );
  AOI22_X1 R2_U880 ( .A1(R2_n2360), .A2(R2_n1271), .B1(R2_n2363), .B2(
        R2_U16_DATA1_13), .ZN(R2_n2185) );
  INV_X1 R2_U879 ( .A(R2_n2185), .ZN(R2_n144) );
  AOI22_X1 R2_U878 ( .A1(R2_n2360), .A2(R2_n1272), .B1(R2_n2363), .B2(
        R2_U16_DATA1_14), .ZN(R2_n2184) );
  INV_X1 R2_U877 ( .A(R2_n2184), .ZN(R2_n145) );
  AOI22_X1 R2_U876 ( .A1(R2_n2360), .A2(R2_n1273), .B1(R2_n2363), .B2(
        R2_U16_DATA1_15), .ZN(R2_n2183) );
  INV_X1 R2_U875 ( .A(R2_n2183), .ZN(R2_n146) );
  AOI22_X1 R2_U874 ( .A1(R2_n2360), .A2(R2_n1274), .B1(R2_n2363), .B2(
        R2_U16_DATA1_16), .ZN(R2_n2182) );
  INV_X1 R2_U873 ( .A(R2_n2182), .ZN(R2_n147) );
  AOI22_X1 R2_U872 ( .A1(R2_n2360), .A2(R2_n1275), .B1(R2_n2362), .B2(
        R2_U16_DATA1_17), .ZN(R2_n2181) );
  INV_X1 R2_U871 ( .A(R2_n2181), .ZN(R2_n148) );
  AOI22_X1 R2_U870 ( .A1(R2_n2360), .A2(R2_n1276), .B1(R2_n2363), .B2(
        R2_U16_DATA1_18), .ZN(R2_n2180) );
  INV_X1 R2_U869 ( .A(R2_n2180), .ZN(R2_n149) );
  AOI22_X1 R2_U868 ( .A1(R2_n2360), .A2(R2_n1277), .B1(R2_n2362), .B2(
        R2_U16_DATA1_19), .ZN(R2_n2179) );
  INV_X1 R2_U867 ( .A(R2_n2179), .ZN(R2_n150) );
  AOI22_X1 R2_U866 ( .A1(R2_n2355), .A2(R2_n1278), .B1(R2_n2362), .B2(
        R2_U16_DATA1_20), .ZN(R2_n2178) );
  INV_X1 R2_U865 ( .A(R2_n2178), .ZN(R2_n151) );
  AOI22_X1 R2_U864 ( .A1(R2_n2360), .A2(R2_n1279), .B1(R2_n2362), .B2(
        R2_U16_DATA1_21), .ZN(R2_n2177) );
  INV_X1 R2_U863 ( .A(R2_n2177), .ZN(R2_n152) );
  AOI22_X1 R2_U862 ( .A1(R2_n2360), .A2(R2_n1280), .B1(R2_n2362), .B2(
        R2_U16_DATA1_22), .ZN(R2_n2176) );
  INV_X1 R2_U861 ( .A(R2_n2176), .ZN(R2_n153) );
  AOI22_X1 R2_U860 ( .A1(R2_n482), .A2(R2_n2350), .B1(R2_n1516), .B2(R2_n2349), 
        .ZN(R2_n2327) );
  INV_X1 R2_U859 ( .A(R2_n2327), .ZN(R2_n2) );
  AOI22_X1 R2_U858 ( .A1(R2_n483), .A2(R2_n2343), .B1(R2_n1517), .B2(R2_n2347), 
        .ZN(R2_n2326) );
  INV_X1 R2_U857 ( .A(R2_n2326), .ZN(R2_n3) );
  AOI22_X1 R2_U856 ( .A1(R2_n484), .A2(R2_n2343), .B1(R2_n1518), .B2(R2_n2348), 
        .ZN(R2_n2325) );
  INV_X1 R2_U855 ( .A(R2_n2325), .ZN(R2_n4) );
  AOI22_X1 R2_U854 ( .A1(R2_n485), .A2(R2_n2343), .B1(R2_n1519), .B2(R2_n2344), 
        .ZN(R2_n2324) );
  INV_X1 R2_U853 ( .A(R2_n2324), .ZN(R2_n5) );
  AOI22_X1 R2_U852 ( .A1(R2_n486), .A2(R2_n2353), .B1(R2_n1520), .B2(R2_n2344), 
        .ZN(R2_n2323) );
  INV_X1 R2_U851 ( .A(R2_n2323), .ZN(R2_n6) );
  AOI22_X1 R2_U850 ( .A1(R2_n487), .A2(R2_n2350), .B1(R2_n1521), .B2(R2_n2344), 
        .ZN(R2_n2322) );
  INV_X1 R2_U849 ( .A(R2_n2322), .ZN(R2_n7) );
  AOI22_X1 R2_U848 ( .A1(R2_n488), .A2(R2_n2200), .B1(R2_n1522), .B2(R2_n2347), 
        .ZN(R2_n2321) );
  INV_X1 R2_U847 ( .A(R2_n2321), .ZN(R2_n8) );
  AOI22_X1 R2_U846 ( .A1(R2_n489), .A2(R2_n2200), .B1(R2_n1523), .B2(R2_n2345), 
        .ZN(R2_n2320) );
  INV_X1 R2_U845 ( .A(R2_n2320), .ZN(R2_n9) );
  AOI22_X1 R2_U844 ( .A1(R2_n490), .A2(R2_n2353), .B1(R2_n1524), .B2(R2_n2345), 
        .ZN(R2_n2319) );
  INV_X1 R2_U843 ( .A(R2_n2319), .ZN(R2_n10) );
  AOI22_X1 R2_U842 ( .A1(R2_n491), .A2(R2_n2353), .B1(R2_n1525), .B2(R2_n2345), 
        .ZN(R2_n2318) );
  INV_X1 R2_U841 ( .A(R2_n2318), .ZN(R2_n11) );
  AOI22_X1 R2_U840 ( .A1(R2_n492), .A2(R2_n2200), .B1(R2_n1526), .B2(R2_n2346), 
        .ZN(R2_n2317) );
  INV_X1 R2_U839 ( .A(R2_n2317), .ZN(R2_n12) );
  AOI22_X1 R2_U838 ( .A1(R2_n493), .A2(R2_n2353), .B1(R2_n1527), .B2(R2_n2349), 
        .ZN(R2_n2316) );
  INV_X1 R2_U837 ( .A(R2_n2316), .ZN(R2_n13) );
  AOI22_X1 R2_U836 ( .A1(R2_n494), .A2(R2_n2343), .B1(R2_n1528), .B2(R2_n2349), 
        .ZN(R2_n2315) );
  INV_X1 R2_U835 ( .A(R2_n2315), .ZN(R2_n14) );
  AOI22_X1 R2_U834 ( .A1(R2_n495), .A2(R2_n2343), .B1(R2_n1529), .B2(R2_n2347), 
        .ZN(R2_n2314) );
  INV_X1 R2_U833 ( .A(R2_n2314), .ZN(R2_n15) );
  AOI22_X1 R2_U832 ( .A1(R2_n496), .A2(R2_n2351), .B1(R2_n1530), .B2(R2_n2348), 
        .ZN(R2_n2313) );
  INV_X1 R2_U831 ( .A(R2_n2313), .ZN(R2_n16) );
  AOI22_X1 R2_U830 ( .A1(R2_n497), .A2(R2_n2200), .B1(R2_n1531), .B2(R2_n2346), 
        .ZN(R2_n2312) );
  INV_X1 R2_U829 ( .A(R2_n2312), .ZN(R2_n17) );
  AOI22_X1 R2_U828 ( .A1(R2_n498), .A2(R2_n2350), .B1(R2_n1532), .B2(R2_n2344), 
        .ZN(R2_n2311) );
  INV_X1 R2_U827 ( .A(R2_n2311), .ZN(R2_n18) );
  AOI22_X1 R2_U826 ( .A1(R2_n499), .A2(R2_n2351), .B1(R2_n1533), .B2(R2_n2349), 
        .ZN(R2_n2310) );
  INV_X1 R2_U825 ( .A(R2_n2310), .ZN(R2_n19) );
  AOI22_X1 R2_U824 ( .A1(R2_n500), .A2(R2_n2343), .B1(R2_n1534), .B2(R2_n2345), 
        .ZN(R2_n2309) );
  INV_X1 R2_U823 ( .A(R2_n2309), .ZN(R2_n20) );
  AOI22_X1 R2_U822 ( .A1(R2_n501), .A2(R2_n2351), .B1(R2_n1535), .B2(R2_n2346), 
        .ZN(R2_n2308) );
  INV_X1 R2_U821 ( .A(R2_n2308), .ZN(R2_n21) );
  AOI22_X1 R2_U820 ( .A1(R2_n502), .A2(R2_n2350), .B1(R2_n1536), .B2(R2_n2344), 
        .ZN(R2_n2307) );
  INV_X1 R2_U819 ( .A(R2_n2307), .ZN(R2_n22) );
  AOI22_X1 R2_U818 ( .A1(R2_n503), .A2(R2_n2350), .B1(R2_n1537), .B2(R2_n2345), 
        .ZN(R2_n2306) );
  INV_X1 R2_U817 ( .A(R2_n2306), .ZN(R2_n23) );
  AOI22_X1 R2_U816 ( .A1(R2_n504), .A2(R2_n2350), .B1(R2_n1538), .B2(R2_n2346), 
        .ZN(R2_n2305) );
  INV_X1 R2_U815 ( .A(R2_n2305), .ZN(R2_n24) );
  AOI22_X1 R2_U814 ( .A1(R2_n505), .A2(R2_n2350), .B1(R2_n1539), .B2(R2_n2347), 
        .ZN(R2_n2304) );
  INV_X1 R2_U813 ( .A(R2_n2304), .ZN(R2_n25) );
  AOI22_X1 R2_U812 ( .A1(R2_n506), .A2(R2_n2352), .B1(R2_n1540), .B2(R2_n2348), 
        .ZN(R2_n2303) );
  INV_X1 R2_U811 ( .A(R2_n2303), .ZN(R2_n26) );
  AOI22_X1 R2_U810 ( .A1(R2_n507), .A2(R2_n2352), .B1(R2_n1541), .B2(R2_n2346), 
        .ZN(R2_n2302) );
  INV_X1 R2_U809 ( .A(R2_n2302), .ZN(R2_n27) );
  AOI22_X1 R2_U808 ( .A1(R2_n508), .A2(R2_n2352), .B1(R2_n1542), .B2(R2_n2347), 
        .ZN(R2_n2301) );
  INV_X1 R2_U807 ( .A(R2_n2301), .ZN(R2_n28) );
  AOI22_X1 R2_U806 ( .A1(R2_n509), .A2(R2_n2352), .B1(R2_n1543), .B2(R2_n2344), 
        .ZN(R2_n2300) );
  INV_X1 R2_U805 ( .A(R2_n2300), .ZN(R2_n29) );
  AOI22_X1 R2_U804 ( .A1(R2_n510), .A2(R2_n2352), .B1(R2_n1544), .B2(R2_n2349), 
        .ZN(R2_n2299) );
  INV_X1 R2_U803 ( .A(R2_n2299), .ZN(R2_n30) );
  AOI22_X1 R2_U802 ( .A1(R2_n511), .A2(R2_n2352), .B1(R2_n1545), .B2(R2_n2347), 
        .ZN(R2_n2298) );
  INV_X1 R2_U801 ( .A(R2_n2298), .ZN(R2_n31) );
  AOI22_X1 R2_U800 ( .A1(R2_n512), .A2(R2_n2351), .B1(R2_n1546), .B2(R2_n2348), 
        .ZN(R2_n2297) );
  INV_X1 R2_U799 ( .A(R2_n2297), .ZN(R2_n32) );
  AOI22_X1 R2_U798 ( .A1(R2_n513), .A2(R2_n2352), .B1(R2_n1547), .B2(R2_n2345), 
        .ZN(R2_n2296) );
  INV_X1 R2_U797 ( .A(R2_n2296), .ZN(R2_n33) );
  AOI22_X1 R2_U796 ( .A1(R2_n514), .A2(R2_n2353), .B1(R2_n1548), .B2(R2_n2344), 
        .ZN(R2_n2295) );
  INV_X1 R2_U795 ( .A(R2_n2295), .ZN(R2_n34) );
  AOI22_X1 R2_U794 ( .A1(R2_n515), .A2(R2_n2353), .B1(R2_n1549), .B2(R2_n2344), 
        .ZN(R2_n2294) );
  INV_X1 R2_U793 ( .A(R2_n2294), .ZN(R2_n35) );
  AOI22_X1 R2_U792 ( .A1(R2_n516), .A2(R2_n2353), .B1(R2_n1550), .B2(R2_n2344), 
        .ZN(R2_n2293) );
  INV_X1 R2_U791 ( .A(R2_n2293), .ZN(R2_n36) );
  AOI22_X1 R2_U790 ( .A1(R2_n517), .A2(R2_n2351), .B1(R2_n1551), .B2(R2_n2346), 
        .ZN(R2_n2292) );
  INV_X1 R2_U789 ( .A(R2_n2292), .ZN(R2_n37) );
  AOI22_X1 R2_U788 ( .A1(R2_n518), .A2(R2_n2352), .B1(R2_n1552), .B2(R2_n2344), 
        .ZN(R2_n2291) );
  INV_X1 R2_U787 ( .A(R2_n2291), .ZN(R2_n38) );
  AOI22_X1 R2_U786 ( .A1(R2_n519), .A2(R2_n2352), .B1(R2_n1553), .B2(R2_n2345), 
        .ZN(R2_n2290) );
  INV_X1 R2_U785 ( .A(R2_n2290), .ZN(R2_n39) );
  AOI22_X1 R2_U784 ( .A1(R2_n520), .A2(R2_n2352), .B1(R2_n1554), .B2(R2_n2349), 
        .ZN(R2_n2289) );
  INV_X1 R2_U783 ( .A(R2_n2289), .ZN(R2_n40) );
  AOI22_X1 R2_U782 ( .A1(R2_n521), .A2(R2_n2352), .B1(R2_n1555), .B2(R2_n2347), 
        .ZN(R2_n2288) );
  INV_X1 R2_U781 ( .A(R2_n2288), .ZN(R2_n41) );
  AOI22_X1 R2_U780 ( .A1(R2_n522), .A2(R2_n2351), .B1(R2_n1556), .B2(R2_n2346), 
        .ZN(R2_n2287) );
  INV_X1 R2_U779 ( .A(R2_n2287), .ZN(R2_n42) );
  AOI22_X1 R2_U778 ( .A1(R2_n523), .A2(R2_n2351), .B1(R2_n1557), .B2(R2_n2344), 
        .ZN(R2_n2286) );
  INV_X1 R2_U777 ( .A(R2_n2286), .ZN(R2_n43) );
  AOI22_X1 R2_U776 ( .A1(R2_n524), .A2(R2_n2351), .B1(R2_n1558), .B2(R2_n2345), 
        .ZN(R2_n2285) );
  INV_X1 R2_U775 ( .A(R2_n2285), .ZN(R2_n44) );
  AOI22_X1 R2_U774 ( .A1(R2_n525), .A2(R2_n2351), .B1(R2_n1559), .B2(R2_n2345), 
        .ZN(R2_n2284) );
  INV_X1 R2_U773 ( .A(R2_n2284), .ZN(R2_n45) );
  AOI22_X1 R2_U772 ( .A1(R2_n526), .A2(R2_n2343), .B1(R2_n1560), .B2(R2_n2345), 
        .ZN(R2_n2283) );
  INV_X1 R2_U771 ( .A(R2_n2283), .ZN(R2_n46) );
  AOI22_X1 R2_U770 ( .A1(R2_n527), .A2(R2_n2343), .B1(R2_n1561), .B2(R2_n2345), 
        .ZN(R2_n2282) );
  INV_X1 R2_U769 ( .A(R2_n2282), .ZN(R2_n47) );
  AOI22_X1 R2_U768 ( .A1(R2_n528), .A2(R2_n2343), .B1(R2_n1562), .B2(R2_n2345), 
        .ZN(R2_n2281) );
  INV_X1 R2_U767 ( .A(R2_n2281), .ZN(R2_n48) );
  AOI22_X1 R2_U766 ( .A1(R2_n529), .A2(R2_n2343), .B1(R2_n1563), .B2(R2_n2345), 
        .ZN(R2_n2280) );
  INV_X1 R2_U765 ( .A(R2_n2280), .ZN(R2_n49) );
  AOI22_X1 R2_U764 ( .A1(R2_n530), .A2(R2_n2352), .B1(R2_n1564), .B2(R2_n2345), 
        .ZN(R2_n2279) );
  INV_X1 R2_U763 ( .A(R2_n2279), .ZN(R2_n50) );
  AOI22_X1 R2_U762 ( .A1(R2_n531), .A2(R2_n2351), .B1(R2_n1565), .B2(R2_n2345), 
        .ZN(R2_n2278) );
  INV_X1 R2_U761 ( .A(R2_n2278), .ZN(R2_n51) );
  AOI22_X1 R2_U760 ( .A1(R2_n532), .A2(R2_n2200), .B1(R2_n1566), .B2(R2_n2344), 
        .ZN(R2_n2277) );
  INV_X1 R2_U759 ( .A(R2_n2277), .ZN(R2_n52) );
  AOI22_X1 R2_U758 ( .A1(R2_n533), .A2(R2_n2343), .B1(R2_n1567), .B2(R2_n2344), 
        .ZN(R2_n2276) );
  INV_X1 R2_U757 ( .A(R2_n2276), .ZN(R2_n53) );
  AOI22_X1 R2_U756 ( .A1(R2_n534), .A2(R2_n2200), .B1(R2_n1568), .B2(R2_n2344), 
        .ZN(R2_n2275) );
  INV_X1 R2_U755 ( .A(R2_n2275), .ZN(R2_n54) );
  AOI22_X1 R2_U754 ( .A1(R2_n535), .A2(R2_n2353), .B1(R2_n1569), .B2(R2_n2344), 
        .ZN(R2_n2274) );
  INV_X1 R2_U753 ( .A(R2_n2274), .ZN(R2_n55) );
  AOI22_X1 R2_U752 ( .A1(R2_n536), .A2(R2_n2352), .B1(R2_n1570), .B2(R2_n2344), 
        .ZN(R2_n2273) );
  INV_X1 R2_U751 ( .A(R2_n2273), .ZN(R2_n56) );
  AOI22_X1 R2_U750 ( .A1(R2_n537), .A2(R2_n2352), .B1(R2_n1571), .B2(R2_n2344), 
        .ZN(R2_n2272) );
  INV_X1 R2_U749 ( .A(R2_n2272), .ZN(R2_n57) );
  AOI22_X1 R2_U748 ( .A1(R2_n538), .A2(R2_n2343), .B1(R2_n1572), .B2(R2_n2346), 
        .ZN(R2_n2271) );
  INV_X1 R2_U747 ( .A(R2_n2271), .ZN(R2_n58) );
  AOI22_X1 R2_U746 ( .A1(R2_n539), .A2(R2_n2352), .B1(R2_n1573), .B2(R2_n2346), 
        .ZN(R2_n2270) );
  INV_X1 R2_U745 ( .A(R2_n2270), .ZN(R2_n59) );
  AOI22_X1 R2_U744 ( .A1(R2_n540), .A2(R2_n2343), .B1(R2_n1574), .B2(R2_n2346), 
        .ZN(R2_n2269) );
  INV_X1 R2_U743 ( .A(R2_n2269), .ZN(R2_n60) );
  AOI22_X1 R2_U742 ( .A1(R2_n541), .A2(R2_n2353), .B1(R2_n1575), .B2(R2_n2346), 
        .ZN(R2_n2268) );
  INV_X1 R2_U741 ( .A(R2_n2268), .ZN(R2_n61) );
  AOI22_X1 R2_U740 ( .A1(R2_n542), .A2(R2_n2343), .B1(R2_n1576), .B2(R2_n2346), 
        .ZN(R2_n2267) );
  INV_X1 R2_U739 ( .A(R2_n2267), .ZN(R2_n62) );
  AOI22_X1 R2_U738 ( .A1(R2_n543), .A2(R2_n2343), .B1(R2_n1577), .B2(R2_n2346), 
        .ZN(R2_n2266) );
  INV_X1 R2_U737 ( .A(R2_n2266), .ZN(R2_n63) );
  AOI22_X1 R2_U736 ( .A1(R2_n544), .A2(R2_n2343), .B1(R2_n1578), .B2(R2_n2346), 
        .ZN(R2_n2265) );
  INV_X1 R2_U735 ( .A(R2_n2265), .ZN(R2_n64) );
  AOI22_X1 R2_U734 ( .A1(R2_n545), .A2(R2_n2343), .B1(R2_n1579), .B2(R2_n2346), 
        .ZN(R2_n2264) );
  INV_X1 R2_U733 ( .A(R2_n2264), .ZN(R2_n65) );
  AOI22_X1 R2_U732 ( .A1(R2_n546), .A2(R2_n2343), .B1(R2_n1580), .B2(R2_n2346), 
        .ZN(R2_n2263) );
  INV_X1 R2_U731 ( .A(R2_n2263), .ZN(R2_n66) );
  AOI22_X1 R2_U730 ( .A1(R2_n547), .A2(R2_n2343), .B1(R2_n1581), .B2(R2_n2345), 
        .ZN(R2_n2262) );
  INV_X1 R2_U729 ( .A(R2_n2262), .ZN(R2_n67) );
  AOI22_X1 R2_U728 ( .A1(R2_n548), .A2(R2_n2350), .B1(R2_n1582), .B2(R2_n2345), 
        .ZN(R2_n2261) );
  INV_X1 R2_U727 ( .A(R2_n2261), .ZN(R2_n68) );
  AOI22_X1 R2_U726 ( .A1(R2_n549), .A2(R2_n2350), .B1(R2_n1583), .B2(R2_n2345), 
        .ZN(R2_n2260) );
  INV_X1 R2_U725 ( .A(R2_n2260), .ZN(R2_n69) );
  AOI22_X1 R2_U724 ( .A1(R2_n550), .A2(R2_n2352), .B1(R2_n1584), .B2(R2_n2346), 
        .ZN(R2_n2259) );
  INV_X1 R2_U723 ( .A(R2_n2259), .ZN(R2_n70) );
  AOI22_X1 R2_U722 ( .A1(R2_n551), .A2(R2_n2350), .B1(R2_n1585), .B2(R2_n2345), 
        .ZN(R2_n2258) );
  INV_X1 R2_U721 ( .A(R2_n2258), .ZN(R2_n71) );
  AOI22_X1 R2_U720 ( .A1(R2_n552), .A2(R2_n2353), .B1(R2_n1586), .B2(R2_n2347), 
        .ZN(R2_n2257) );
  INV_X1 R2_U719 ( .A(R2_n2257), .ZN(R2_n72) );
  AOI22_X1 R2_U718 ( .A1(R2_n553), .A2(R2_n2353), .B1(R2_n1587), .B2(R2_n2347), 
        .ZN(R2_n2256) );
  INV_X1 R2_U717 ( .A(R2_n2256), .ZN(R2_n73) );
  AOI22_X1 R2_U716 ( .A1(R2_n554), .A2(R2_n2200), .B1(R2_n1588), .B2(R2_n2349), 
        .ZN(R2_n2255) );
  INV_X1 R2_U715 ( .A(R2_n2255), .ZN(R2_n74) );
  AOI22_X1 R2_U714 ( .A1(R2_n555), .A2(R2_n2200), .B1(R2_n1589), .B2(R2_n2347), 
        .ZN(R2_n2254) );
  INV_X1 R2_U713 ( .A(R2_n2254), .ZN(R2_n75) );
  AOI22_X1 R2_U712 ( .A1(R2_n556), .A2(R2_n2353), .B1(R2_n1590), .B2(R2_n2348), 
        .ZN(R2_n2253) );
  INV_X1 R2_U711 ( .A(R2_n2253), .ZN(R2_n76) );
  AOI22_X1 R2_U710 ( .A1(R2_n557), .A2(R2_n2352), .B1(R2_n1591), .B2(R2_n2348), 
        .ZN(R2_n2252) );
  INV_X1 R2_U709 ( .A(R2_n2252), .ZN(R2_n77) );
  AOI22_X1 R2_U708 ( .A1(R2_n558), .A2(R2_n2350), .B1(R2_n1592), .B2(R2_n2344), 
        .ZN(R2_n2251) );
  INV_X1 R2_U707 ( .A(R2_n2251), .ZN(R2_n78) );
  AOI22_X1 R2_U706 ( .A1(R2_n559), .A2(R2_n2350), .B1(R2_n1593), .B2(R2_n2344), 
        .ZN(R2_n2250) );
  INV_X1 R2_U705 ( .A(R2_n2250), .ZN(R2_n79) );
  AOI22_X1 R2_U704 ( .A1(R2_n560), .A2(R2_n2200), .B1(R2_n1594), .B2(R2_n2345), 
        .ZN(R2_n2249) );
  INV_X1 R2_U703 ( .A(R2_n2249), .ZN(R2_n80) );
  AOI22_X1 R2_U702 ( .A1(R2_n561), .A2(R2_n2353), .B1(R2_n1595), .B2(R2_n2346), 
        .ZN(R2_n2248) );
  INV_X1 R2_U701 ( .A(R2_n2248), .ZN(R2_n81) );
  AOI22_X1 R2_U700 ( .A1(R2_n562), .A2(R2_n2350), .B1(R2_n1596), .B2(R2_n2344), 
        .ZN(R2_n2247) );
  INV_X1 R2_U699 ( .A(R2_n2247), .ZN(R2_n82) );
  AOI22_X1 R2_U698 ( .A1(R2_n563), .A2(R2_n2200), .B1(R2_n1597), .B2(R2_n2349), 
        .ZN(R2_n2246) );
  INV_X1 R2_U697 ( .A(R2_n2246), .ZN(R2_n83) );
  AOI22_X1 R2_U696 ( .A1(R2_n564), .A2(R2_n2352), .B1(R2_n1598), .B2(R2_n2349), 
        .ZN(R2_n2245) );
  INV_X1 R2_U695 ( .A(R2_n2245), .ZN(R2_n84) );
  AOI22_X1 R2_U694 ( .A1(R2_n565), .A2(R2_n2353), .B1(R2_n1599), .B2(R2_n2349), 
        .ZN(R2_n2244) );
  INV_X1 R2_U693 ( .A(R2_n2244), .ZN(R2_n85) );
  AOI22_X1 R2_U692 ( .A1(R2_n566), .A2(R2_n2200), .B1(R2_n1600), .B2(R2_n2345), 
        .ZN(R2_n2243) );
  INV_X1 R2_U691 ( .A(R2_n2243), .ZN(R2_n86) );
  AOI22_X1 R2_U690 ( .A1(R2_n567), .A2(R2_n2353), .B1(R2_n1601), .B2(R2_n2349), 
        .ZN(R2_n2242) );
  INV_X1 R2_U689 ( .A(R2_n2242), .ZN(R2_n87) );
  AOI22_X1 R2_U688 ( .A1(R2_n568), .A2(R2_n2350), .B1(R2_n1602), .B2(R2_n2349), 
        .ZN(R2_n2241) );
  INV_X1 R2_U687 ( .A(R2_n2241), .ZN(R2_n88) );
  AOI22_X1 R2_U686 ( .A1(R2_n569), .A2(R2_n2200), .B1(R2_n1603), .B2(R2_n2349), 
        .ZN(R2_n2240) );
  INV_X1 R2_U685 ( .A(R2_n2240), .ZN(R2_n89) );
  AOI22_X1 R2_U684 ( .A1(R2_n570), .A2(R2_n2350), .B1(R2_n1604), .B2(R2_n2349), 
        .ZN(R2_n2239) );
  INV_X1 R2_U683 ( .A(R2_n2239), .ZN(R2_n90) );
  AOI22_X1 R2_U682 ( .A1(R2_n571), .A2(R2_n2350), .B1(R2_n1605), .B2(R2_n2348), 
        .ZN(R2_n2238) );
  INV_X1 R2_U681 ( .A(R2_n2238), .ZN(R2_n91) );
  AOI22_X1 R2_U680 ( .A1(R2_n572), .A2(R2_n2350), .B1(R2_n1606), .B2(R2_n2349), 
        .ZN(R2_n2237) );
  INV_X1 R2_U679 ( .A(R2_n2237), .ZN(R2_n92) );
  AOI22_X1 R2_U678 ( .A1(R2_n573), .A2(R2_n2353), .B1(R2_n1607), .B2(R2_n2349), 
        .ZN(R2_n2236) );
  INV_X1 R2_U677 ( .A(R2_n2236), .ZN(R2_n93) );
  AOI22_X1 R2_U676 ( .A1(R2_n574), .A2(R2_n2200), .B1(R2_n1608), .B2(R2_n2349), 
        .ZN(R2_n2235) );
  INV_X1 R2_U675 ( .A(R2_n2235), .ZN(R2_n94) );
  AOI22_X1 R2_U674 ( .A1(R2_n575), .A2(R2_n2350), .B1(R2_n1609), .B2(R2_n2344), 
        .ZN(R2_n2234) );
  INV_X1 R2_U673 ( .A(R2_n2234), .ZN(R2_n95) );
  AOI22_X1 R2_U672 ( .A1(R2_n576), .A2(R2_n2353), .B1(R2_n1610), .B2(R2_n2349), 
        .ZN(R2_n2233) );
  INV_X1 R2_U671 ( .A(R2_n2233), .ZN(R2_n96) );
  AOI22_X1 R2_U670 ( .A1(R2_n577), .A2(R2_n2350), .B1(R2_n1611), .B2(R2_n2345), 
        .ZN(R2_n2232) );
  INV_X1 R2_U669 ( .A(R2_n2232), .ZN(R2_n97) );
  AOI22_X1 R2_U668 ( .A1(R2_n578), .A2(R2_n2200), .B1(R2_n1612), .B2(R2_n2347), 
        .ZN(R2_n2231) );
  INV_X1 R2_U667 ( .A(R2_n2231), .ZN(R2_n98) );
  AOI22_X1 R2_U666 ( .A1(R2_n579), .A2(R2_n2200), .B1(R2_n1613), .B2(R2_n2346), 
        .ZN(R2_n2230) );
  INV_X1 R2_U665 ( .A(R2_n2230), .ZN(R2_n99) );
  AOI22_X1 R2_U664 ( .A1(R2_n580), .A2(R2_n2353), .B1(R2_n1614), .B2(R2_n2347), 
        .ZN(R2_n2229) );
  INV_X1 R2_U663 ( .A(R2_n2229), .ZN(R2_n100) );
  AOI22_X1 R2_U662 ( .A1(R2_n581), .A2(R2_n2351), .B1(R2_n1615), .B2(R2_n2348), 
        .ZN(R2_n2228) );
  INV_X1 R2_U661 ( .A(R2_n2228), .ZN(R2_n101) );
  AOI22_X1 R2_U660 ( .A1(R2_n582), .A2(R2_n2352), .B1(R2_n1616), .B2(R2_n2349), 
        .ZN(R2_n2227) );
  INV_X1 R2_U659 ( .A(R2_n2227), .ZN(R2_n102) );
  AOI22_X1 R2_U658 ( .A1(R2_n583), .A2(R2_n2350), .B1(R2_n1617), .B2(R2_n2344), 
        .ZN(R2_n2226) );
  INV_X1 R2_U657 ( .A(R2_n2226), .ZN(R2_n103) );
  AOI22_X1 R2_U656 ( .A1(R2_n584), .A2(R2_n2351), .B1(R2_n1618), .B2(R2_n2345), 
        .ZN(R2_n2225) );
  INV_X1 R2_U655 ( .A(R2_n2225), .ZN(R2_n104) );
  AOI22_X1 R2_U654 ( .A1(R2_n585), .A2(R2_n2351), .B1(R2_n1619), .B2(R2_n2349), 
        .ZN(R2_n2224) );
  INV_X1 R2_U653 ( .A(R2_n2224), .ZN(R2_n105) );
  AOI22_X1 R2_U652 ( .A1(R2_n586), .A2(R2_n2350), .B1(R2_n1620), .B2(R2_n2347), 
        .ZN(R2_n2223) );
  INV_X1 R2_U651 ( .A(R2_n2223), .ZN(R2_n106) );
  AOI22_X1 R2_U650 ( .A1(R2_n587), .A2(R2_n2352), .B1(R2_n1621), .B2(R2_n2347), 
        .ZN(R2_n2222) );
  INV_X1 R2_U649 ( .A(R2_n2222), .ZN(R2_n107) );
  AOI22_X1 R2_U648 ( .A1(R2_n588), .A2(R2_n2351), .B1(R2_n1622), .B2(R2_n2347), 
        .ZN(R2_n2221) );
  INV_X1 R2_U647 ( .A(R2_n2221), .ZN(R2_n108) );
  AOI22_X1 R2_U646 ( .A1(R2_n589), .A2(R2_n2350), .B1(R2_n1623), .B2(R2_n2347), 
        .ZN(R2_n2220) );
  INV_X1 R2_U645 ( .A(R2_n2220), .ZN(R2_n109) );
  AOI22_X1 R2_U644 ( .A1(R2_n590), .A2(R2_n2200), .B1(R2_n1624), .B2(R2_n2347), 
        .ZN(R2_n2219) );
  INV_X1 R2_U643 ( .A(R2_n2219), .ZN(R2_n110) );
  AOI22_X1 R2_U642 ( .A1(R2_n591), .A2(R2_n2351), .B1(R2_n1625), .B2(R2_n2347), 
        .ZN(R2_n2218) );
  INV_X1 R2_U641 ( .A(R2_n2218), .ZN(R2_n111) );
  AOI22_X1 R2_U640 ( .A1(R2_n592), .A2(R2_n2352), .B1(R2_n1626), .B2(R2_n2347), 
        .ZN(R2_n2217) );
  INV_X1 R2_U639 ( .A(R2_n2217), .ZN(R2_n112) );
  AOI22_X1 R2_U638 ( .A1(R2_n593), .A2(R2_n2352), .B1(R2_n1627), .B2(R2_n2347), 
        .ZN(R2_n2216) );
  INV_X1 R2_U637 ( .A(R2_n2216), .ZN(R2_n113) );
  AOI22_X1 R2_U636 ( .A1(R2_n594), .A2(R2_n2200), .B1(R2_n1628), .B2(R2_n2347), 
        .ZN(R2_n2215) );
  INV_X1 R2_U635 ( .A(R2_n2215), .ZN(R2_n114) );
  AOI22_X1 R2_U634 ( .A1(R2_n595), .A2(R2_n2200), .B1(R2_n1629), .B2(R2_n2348), 
        .ZN(R2_n2214) );
  INV_X1 R2_U633 ( .A(R2_n2214), .ZN(R2_n115) );
  AOI22_X1 R2_U632 ( .A1(R2_n596), .A2(R2_n2353), .B1(R2_n1630), .B2(R2_n2344), 
        .ZN(R2_n2213) );
  INV_X1 R2_U631 ( .A(R2_n2213), .ZN(R2_n116) );
  AOI22_X1 R2_U630 ( .A1(R2_n597), .A2(R2_n2200), .B1(R2_n1631), .B2(R2_n2346), 
        .ZN(R2_n2212) );
  INV_X1 R2_U629 ( .A(R2_n2212), .ZN(R2_n117) );
  AOI22_X1 R2_U628 ( .A1(R2_n598), .A2(R2_n2353), .B1(R2_n1632), .B2(R2_n2348), 
        .ZN(R2_n2211) );
  INV_X1 R2_U627 ( .A(R2_n2211), .ZN(R2_n118) );
  AOI22_X1 R2_U626 ( .A1(R2_n599), .A2(R2_n2353), .B1(R2_n1633), .B2(R2_n2349), 
        .ZN(R2_n2210) );
  INV_X1 R2_U625 ( .A(R2_n2210), .ZN(R2_n119) );
  AOI22_X1 R2_U624 ( .A1(R2_n600), .A2(R2_n2350), .B1(R2_n1634), .B2(R2_n2349), 
        .ZN(R2_n2209) );
  INV_X1 R2_U623 ( .A(R2_n2209), .ZN(R2_n120) );
  AOI22_X1 R2_U622 ( .A1(R2_n601), .A2(R2_n2353), .B1(R2_n1635), .B2(R2_n2348), 
        .ZN(R2_n2208) );
  INV_X1 R2_U621 ( .A(R2_n2208), .ZN(R2_n121) );
  AOI22_X1 R2_U620 ( .A1(R2_n602), .A2(R2_n2353), .B1(R2_n1636), .B2(R2_n2347), 
        .ZN(R2_n2207) );
  INV_X1 R2_U619 ( .A(R2_n2207), .ZN(R2_n122) );
  AOI22_X1 R2_U618 ( .A1(R2_n603), .A2(R2_n2351), .B1(R2_n1637), .B2(R2_n2348), 
        .ZN(R2_n2206) );
  INV_X1 R2_U617 ( .A(R2_n2206), .ZN(R2_n123) );
  AOI22_X1 R2_U616 ( .A1(R2_n604), .A2(R2_n2353), .B1(R2_n1638), .B2(R2_n2348), 
        .ZN(R2_n2205) );
  INV_X1 R2_U615 ( .A(R2_n2205), .ZN(R2_n124) );
  AOI22_X1 R2_U614 ( .A1(R2_n605), .A2(R2_n2351), .B1(R2_n1639), .B2(R2_n2348), 
        .ZN(R2_n2204) );
  INV_X1 R2_U613 ( .A(R2_n2204), .ZN(R2_n125) );
  AOI22_X1 R2_U612 ( .A1(R2_n606), .A2(R2_n2353), .B1(R2_n1640), .B2(R2_n2348), 
        .ZN(R2_n2203) );
  INV_X1 R2_U611 ( .A(R2_n2203), .ZN(R2_n126) );
  AOI22_X1 R2_U610 ( .A1(R2_n607), .A2(R2_n2200), .B1(R2_n1641), .B2(R2_n2348), 
        .ZN(R2_n2202) );
  INV_X1 R2_U609 ( .A(R2_n2202), .ZN(R2_n127) );
  AOI22_X1 R2_U608 ( .A1(R2_n608), .A2(R2_n2353), .B1(R2_n1642), .B2(R2_n2348), 
        .ZN(R2_n2201) );
  INV_X1 R2_U607 ( .A(R2_n2201), .ZN(R2_n128) );
  AOI22_X1 R2_U606 ( .A1(R2_n609), .A2(R2_n2353), .B1(R2_n1643), .B2(R2_n2348), 
        .ZN(R2_n2199) );
  INV_X1 R2_U605 ( .A(R2_n2199), .ZN(R2_n129) );
  AOI22_X1 R2_U604 ( .A1(n3263), .A2(R2_n2384), .B1(R2_n[616]), .B2(R2_n2379), 
        .ZN(R2_n1938) );
  INV_X1 R2_U603 ( .A(R2_n1938), .ZN(R2_n1030) );
  AOI22_X1 R2_U602 ( .A1(n3264), .A2(R2_n2385), .B1(R2_n[617]), .B2(R2_n2378), 
        .ZN(R2_n1937) );
  INV_X1 R2_U601 ( .A(R2_n1937), .ZN(R2_n1031) );
  AOI22_X1 R2_U600 ( .A1(n3265), .A2(R2_n2383), .B1(R2_n[618]), .B2(R2_n2378), 
        .ZN(R2_n1936) );
  INV_X1 R2_U599 ( .A(R2_n1936), .ZN(R2_n1032) );
  AOI22_X1 R2_U598 ( .A1(n3266), .A2(R2_n2375), .B1(R2_n[619]), .B2(R2_n2381), 
        .ZN(R2_n1935) );
  INV_X1 R2_U597 ( .A(R2_n1935), .ZN(R2_n1033) );
  AOI22_X1 R2_U596 ( .A1(n3267), .A2(R2_n2383), .B1(R2_n[620]), .B2(R2_n2378), 
        .ZN(R2_n1934) );
  INV_X1 R2_U595 ( .A(R2_n1934), .ZN(R2_n1034) );
  AOI22_X1 R2_U594 ( .A1(n3268), .A2(R2_n2383), .B1(R2_n[621]), .B2(R2_n2382), 
        .ZN(R2_n1933) );
  INV_X1 R2_U593 ( .A(R2_n1933), .ZN(R2_n1035) );
  AOI22_X1 R2_U592 ( .A1(n3269), .A2(R2_n2375), .B1(R2_n[622]), .B2(R2_n2381), 
        .ZN(R2_n1932) );
  INV_X1 R2_U591 ( .A(R2_n1932), .ZN(R2_n1036) );
  AOI22_X1 R2_U590 ( .A1(n3270), .A2(R2_n2385), .B1(R2_n[623]), .B2(R2_n2378), 
        .ZN(R2_n1931) );
  INV_X1 R2_U589 ( .A(R2_n1931), .ZN(R2_n1037) );
  AOI22_X1 R2_U588 ( .A1(n3271), .A2(R2_n2376), .B1(R2_n[624]), .B2(R2_n2378), 
        .ZN(R2_n1930) );
  INV_X1 R2_U587 ( .A(R2_n1930), .ZN(R2_n1038) );
  AOI22_X1 R2_U586 ( .A1(n3272), .A2(R2_n2376), .B1(R2_n[625]), .B2(R2_n2379), 
        .ZN(R2_n1929) );
  INV_X1 R2_U585 ( .A(R2_n1929), .ZN(R2_n1039) );
  AOI22_X1 R2_U584 ( .A1(n3273), .A2(R2_n2376), .B1(R2_n[626]), .B2(R2_n2378), 
        .ZN(R2_n1928) );
  INV_X1 R2_U583 ( .A(R2_n1928), .ZN(R2_n1040) );
  AOI22_X1 R2_U582 ( .A1(n3274), .A2(R2_n2375), .B1(R2_n[627]), .B2(R2_n2377), 
        .ZN(R2_n1927) );
  INV_X1 R2_U581 ( .A(R2_n1927), .ZN(R2_n1041) );
  AOI22_X1 R2_U580 ( .A1(n3275), .A2(R2_n2376), .B1(R2_n[628]), .B2(R2_n2378), 
        .ZN(R2_n1926) );
  INV_X1 R2_U579 ( .A(R2_n1926), .ZN(R2_n1042) );
  AOI22_X1 R2_U578 ( .A1(n3276), .A2(R2_n1811), .B1(R2_n[629]), .B2(R2_n2377), 
        .ZN(R2_n1925) );
  INV_X1 R2_U577 ( .A(R2_n1925), .ZN(R2_n1043) );
  AOI22_X1 R2_U576 ( .A1(n3277), .A2(R2_n2384), .B1(R2_n[630]), .B2(R2_n2382), 
        .ZN(R2_n1924) );
  INV_X1 R2_U575 ( .A(R2_n1924), .ZN(R2_n1044) );
  AOI22_X1 R2_U574 ( .A1(n3278), .A2(R2_n2385), .B1(R2_n[631]), .B2(R2_n2381), 
        .ZN(R2_n1923) );
  INV_X1 R2_U573 ( .A(R2_n1923), .ZN(R2_n1045) );
  AOI22_X1 R2_U572 ( .A1(n3279), .A2(R2_n1811), .B1(R2_n[632]), .B2(R2_n2377), 
        .ZN(R2_n1922) );
  INV_X1 R2_U571 ( .A(R2_n1922), .ZN(R2_n1046) );
  AOI22_X1 R2_U570 ( .A1(n3280), .A2(R2_n2375), .B1(R2_n[633]), .B2(R2_n2380), 
        .ZN(R2_n1921) );
  INV_X1 R2_U569 ( .A(R2_n1921), .ZN(R2_n1047) );
  AOI22_X1 R2_U568 ( .A1(n3281), .A2(R2_n2376), .B1(R2_n[634]), .B2(R2_n2378), 
        .ZN(R2_n1920) );
  INV_X1 R2_U567 ( .A(R2_n1920), .ZN(R2_n1048) );
  AOI22_X1 R2_U566 ( .A1(n3282), .A2(R2_n1811), .B1(R2_n[635]), .B2(R2_n2379), 
        .ZN(R2_n1919) );
  INV_X1 R2_U565 ( .A(R2_n1919), .ZN(R2_n1049) );
  AOI22_X1 R2_U564 ( .A1(n3283), .A2(R2_n2385), .B1(R2_n[636]), .B2(R2_n2379), 
        .ZN(R2_n1918) );
  INV_X1 R2_U563 ( .A(R2_n1918), .ZN(R2_n1050) );
  AOI22_X1 R2_U562 ( .A1(n3284), .A2(R2_n2385), .B1(R2_n[637]), .B2(R2_n2377), 
        .ZN(R2_n1917) );
  INV_X1 R2_U561 ( .A(R2_n1917), .ZN(R2_n1051) );
  AOI22_X1 R2_U560 ( .A1(n3285), .A2(R2_n2385), .B1(R2_n[638]), .B2(R2_n2380), 
        .ZN(R2_n1916) );
  INV_X1 R2_U559 ( .A(R2_n1916), .ZN(R2_n1052) );
  AOI22_X1 R2_U558 ( .A1(n3286), .A2(R2_n2385), .B1(R2_n[639]), .B2(R2_n2379), 
        .ZN(R2_n1915) );
  INV_X1 R2_U557 ( .A(R2_n1915), .ZN(R2_n1053) );
  AOI22_X1 R2_U556 ( .A1(n3287), .A2(R2_n2384), .B1(R2_n[640]), .B2(R2_n2379), 
        .ZN(R2_n1914) );
  INV_X1 R2_U555 ( .A(R2_n1914), .ZN(R2_n1054) );
  AOI22_X1 R2_U554 ( .A1(n3288), .A2(R2_n2384), .B1(R2_n[641]), .B2(R2_n2382), 
        .ZN(R2_n1913) );
  INV_X1 R2_U553 ( .A(R2_n1913), .ZN(R2_n1055) );
  AOI22_X1 R2_U552 ( .A1(n3289), .A2(R2_n2384), .B1(R2_n[642]), .B2(R2_n2381), 
        .ZN(R2_n1912) );
  INV_X1 R2_U551 ( .A(R2_n1912), .ZN(R2_n1056) );
  AOI22_X1 R2_U550 ( .A1(n3290), .A2(R2_n2384), .B1(R2_n[643]), .B2(R2_n2379), 
        .ZN(R2_n1911) );
  INV_X1 R2_U549 ( .A(R2_n1911), .ZN(R2_n1057) );
  AOI22_X1 R2_U548 ( .A1(n3291), .A2(R2_n2383), .B1(R2_n[644]), .B2(R2_n2378), 
        .ZN(R2_n1910) );
  INV_X1 R2_U547 ( .A(R2_n1910), .ZN(R2_n1058) );
  AOI22_X1 R2_U546 ( .A1(n3292), .A2(R2_n2383), .B1(R2_n[645]), .B2(R2_n2382), 
        .ZN(R2_n1909) );
  INV_X1 R2_U545 ( .A(R2_n1909), .ZN(R2_n1059) );
  AOI22_X1 R2_U544 ( .A1(n3293), .A2(R2_n2383), .B1(R2_n[646]), .B2(R2_n2381), 
        .ZN(R2_n1908) );
  INV_X1 R2_U543 ( .A(R2_n1908), .ZN(R2_n1060) );
  AOI22_X1 R2_U542 ( .A1(n3294), .A2(R2_n2383), .B1(R2_n[647]), .B2(R2_n2377), 
        .ZN(R2_n1907) );
  INV_X1 R2_U541 ( .A(R2_n1907), .ZN(R2_n1061) );
  AOI22_X1 R2_U540 ( .A1(n3295), .A2(R2_n2384), .B1(R2_n[648]), .B2(R2_n2380), 
        .ZN(R2_n1906) );
  INV_X1 R2_U539 ( .A(R2_n1906), .ZN(R2_n1062) );
  AOI22_X1 R2_U538 ( .A1(n3296), .A2(R2_n2376), .B1(R2_n[649]), .B2(R2_n2379), 
        .ZN(R2_n1905) );
  INV_X1 R2_U537 ( .A(R2_n1905), .ZN(R2_n1063) );
  AOI22_X1 R2_U536 ( .A1(n3297), .A2(R2_n2376), .B1(R2_n[650]), .B2(R2_n2378), 
        .ZN(R2_n1904) );
  INV_X1 R2_U535 ( .A(R2_n1904), .ZN(R2_n1064) );
  AOI22_X1 R2_U534 ( .A1(n3298), .A2(R2_n2385), .B1(R2_n[651]), .B2(R2_n2382), 
        .ZN(R2_n1903) );
  INV_X1 R2_U533 ( .A(R2_n1903), .ZN(R2_n1065) );
  AOI22_X1 R2_U532 ( .A1(n3299), .A2(R2_n1811), .B1(R2_n[652]), .B2(R2_n2379), 
        .ZN(R2_n1902) );
  INV_X1 R2_U531 ( .A(R2_n1902), .ZN(R2_n1066) );
  AOI22_X1 R2_U530 ( .A1(n3300), .A2(R2_n1811), .B1(R2_n[653]), .B2(R2_n2377), 
        .ZN(R2_n1901) );
  INV_X1 R2_U529 ( .A(R2_n1901), .ZN(R2_n1067) );
  AOI22_X1 R2_U528 ( .A1(n3301), .A2(R2_n1811), .B1(R2_n[654]), .B2(R2_n2382), 
        .ZN(R2_n1900) );
  INV_X1 R2_U527 ( .A(R2_n1900), .ZN(R2_n1068) );
  AOI22_X1 R2_U526 ( .A1(n3302), .A2(R2_n1811), .B1(R2_n[655]), .B2(R2_n2377), 
        .ZN(R2_n1899) );
  INV_X1 R2_U525 ( .A(R2_n1899), .ZN(R2_n1069) );
  AOI22_X1 R2_U524 ( .A1(n3303), .A2(R2_n2384), .B1(R2_n[656]), .B2(R2_n2380), 
        .ZN(R2_n1898) );
  INV_X1 R2_U523 ( .A(R2_n1898), .ZN(R2_n1070) );
  AOI22_X1 R2_U522 ( .A1(n3304), .A2(R2_n2385), .B1(R2_n[657]), .B2(R2_n2380), 
        .ZN(R2_n1897) );
  INV_X1 R2_U521 ( .A(R2_n1897), .ZN(R2_n1071) );
  AOI22_X1 R2_U520 ( .A1(n3305), .A2(R2_n2383), .B1(R2_n[658]), .B2(R2_n2381), 
        .ZN(R2_n1896) );
  INV_X1 R2_U519 ( .A(R2_n1896), .ZN(R2_n1072) );
  AOI22_X1 R2_U518 ( .A1(n3306), .A2(R2_n2383), .B1(R2_n[659]), .B2(R2_n2377), 
        .ZN(R2_n1895) );
  INV_X1 R2_U517 ( .A(R2_n1895), .ZN(R2_n1073) );
  AOI22_X1 R2_U516 ( .A1(n3307), .A2(R2_n1811), .B1(R2_n[660]), .B2(R2_n2380), 
        .ZN(R2_n1894) );
  INV_X1 R2_U515 ( .A(R2_n1894), .ZN(R2_n1074) );
  AOI22_X1 R2_U514 ( .A1(n3308), .A2(R2_n1811), .B1(R2_n[661]), .B2(R2_n2378), 
        .ZN(R2_n1893) );
  INV_X1 R2_U513 ( .A(R2_n1893), .ZN(R2_n1075) );
  AOI22_X1 R2_U512 ( .A1(n3309), .A2(R2_n1811), .B1(R2_n[662]), .B2(R2_n2379), 
        .ZN(R2_n1892) );
  INV_X1 R2_U511 ( .A(R2_n1892), .ZN(R2_n1076) );
  AOI22_X1 R2_U510 ( .A1(n3310), .A2(R2_n1811), .B1(R2_n[663]), .B2(R2_n2380), 
        .ZN(R2_n1891) );
  INV_X1 R2_U509 ( .A(R2_n1891), .ZN(R2_n1077) );
  AOI22_X1 R2_U508 ( .A1(n3311), .A2(R2_n2376), .B1(R2_n[664]), .B2(R2_n2382), 
        .ZN(R2_n1890) );
  INV_X1 R2_U507 ( .A(R2_n1890), .ZN(R2_n1078) );
  AOI22_X1 R2_U506 ( .A1(n3312), .A2(R2_n2376), .B1(R2_n[665]), .B2(R2_n2381), 
        .ZN(R2_n1889) );
  INV_X1 R2_U505 ( .A(R2_n1889), .ZN(R2_n1079) );
  AOI22_X1 R2_U504 ( .A1(n3313), .A2(R2_n2376), .B1(R2_n[666]), .B2(R2_n2377), 
        .ZN(R2_n1888) );
  INV_X1 R2_U503 ( .A(R2_n1888), .ZN(R2_n1080) );
  AOI22_X1 R2_U502 ( .A1(n3314), .A2(R2_n2376), .B1(R2_n[667]), .B2(R2_n2377), 
        .ZN(R2_n1887) );
  INV_X1 R2_U501 ( .A(R2_n1887), .ZN(R2_n1081) );
  AOI22_X1 R2_U500 ( .A1(n3315), .A2(R2_n2385), .B1(R2_n[668]), .B2(R2_n2380), 
        .ZN(R2_n1886) );
  INV_X1 R2_U499 ( .A(R2_n1886), .ZN(R2_n1082) );
  AOI22_X1 R2_U498 ( .A1(n3316), .A2(R2_n2384), .B1(R2_n[669]), .B2(R2_n2380), 
        .ZN(R2_n1885) );
  INV_X1 R2_U497 ( .A(R2_n1885), .ZN(R2_n1083) );
  AOI22_X1 R2_U496 ( .A1(n3317), .A2(R2_n2383), .B1(R2_n[670]), .B2(R2_n2380), 
        .ZN(R2_n1884) );
  INV_X1 R2_U495 ( .A(R2_n1884), .ZN(R2_n1084) );
  AOI22_X1 R2_U494 ( .A1(n3318), .A2(R2_n2384), .B1(R2_n[671]), .B2(R2_n2378), 
        .ZN(R2_n1883) );
  INV_X1 R2_U493 ( .A(R2_n1883), .ZN(R2_n1085) );
  AOI22_X1 R2_U492 ( .A1(n3319), .A2(R2_n2383), .B1(R2_n[672]), .B2(R2_n2382), 
        .ZN(R2_n1882) );
  INV_X1 R2_U491 ( .A(R2_n1882), .ZN(R2_n1086) );
  AOI22_X1 R2_U490 ( .A1(n3320), .A2(R2_n1811), .B1(R2_n[673]), .B2(R2_n2382), 
        .ZN(R2_n1881) );
  INV_X1 R2_U489 ( .A(R2_n1881), .ZN(R2_n1087) );
  AOI22_X1 R2_U488 ( .A1(n3321), .A2(R2_n2375), .B1(R2_n[674]), .B2(R2_n2381), 
        .ZN(R2_n1880) );
  INV_X1 R2_U487 ( .A(R2_n1880), .ZN(R2_n1088) );
  AOI22_X1 R2_U486 ( .A1(n3322), .A2(R2_n1811), .B1(R2_n[675]), .B2(R2_n2377), 
        .ZN(R2_n1879) );
  INV_X1 R2_U485 ( .A(R2_n1879), .ZN(R2_n1089) );
  AOI22_X1 R2_U484 ( .A1(n3323), .A2(R2_n2385), .B1(R2_n[676]), .B2(R2_n2380), 
        .ZN(R2_n1878) );
  INV_X1 R2_U483 ( .A(R2_n1878), .ZN(R2_n1090) );
  AOI22_X1 R2_U482 ( .A1(n3324), .A2(R2_n1811), .B1(R2_n[677]), .B2(R2_n2379), 
        .ZN(R2_n1877) );
  INV_X1 R2_U481 ( .A(R2_n1877), .ZN(R2_n1091) );
  AOI22_X1 R2_U480 ( .A1(n3325), .A2(R2_n2375), .B1(R2_n[678]), .B2(R2_n2381), 
        .ZN(R2_n1876) );
  INV_X1 R2_U479 ( .A(R2_n1876), .ZN(R2_n1092) );
  AOI22_X1 R2_U478 ( .A1(n3326), .A2(R2_n2376), .B1(R2_n[679]), .B2(R2_n2377), 
        .ZN(R2_n1875) );
  INV_X1 R2_U477 ( .A(R2_n1875), .ZN(R2_n1093) );
  AOI22_X1 R2_U476 ( .A1(n3327), .A2(R2_n2383), .B1(R2_n[680]), .B2(R2_n2377), 
        .ZN(R2_n1874) );
  INV_X1 R2_U475 ( .A(R2_n1874), .ZN(R2_n1094) );
  AOI22_X1 R2_U474 ( .A1(n3328), .A2(R2_n2376), .B1(R2_n[681]), .B2(R2_n2377), 
        .ZN(R2_n1873) );
  INV_X1 R2_U473 ( .A(R2_n1873), .ZN(R2_n1095) );
  AOI22_X1 R2_U472 ( .A1(n3329), .A2(R2_n2376), .B1(R2_n[682]), .B2(R2_n2377), 
        .ZN(R2_n1872) );
  INV_X1 R2_U471 ( .A(R2_n1872), .ZN(R2_n1096) );
  AOI22_X1 R2_U470 ( .A1(n3330), .A2(R2_n2384), .B1(R2_n[683]), .B2(R2_n2377), 
        .ZN(R2_n1871) );
  INV_X1 R2_U469 ( .A(R2_n1871), .ZN(R2_n1097) );
  AOI22_X1 R2_U468 ( .A1(n3331), .A2(R2_n2384), .B1(R2_n[684]), .B2(R2_n2377), 
        .ZN(R2_n1870) );
  INV_X1 R2_U467 ( .A(R2_n1870), .ZN(R2_n1098) );
  AOI22_X1 R2_U466 ( .A1(n3332), .A2(R2_n2384), .B1(R2_n[685]), .B2(R2_n2377), 
        .ZN(R2_n1869) );
  INV_X1 R2_U465 ( .A(R2_n1869), .ZN(R2_n1099) );
  AOI22_X1 R2_U464 ( .A1(n3333), .A2(R2_n2376), .B1(R2_n[686]), .B2(R2_n2377), 
        .ZN(R2_n1868) );
  INV_X1 R2_U463 ( .A(R2_n1868), .ZN(R2_n1100) );
  AOI22_X1 R2_U462 ( .A1(n3334), .A2(R2_n2375), .B1(R2_n[687]), .B2(R2_n2377), 
        .ZN(R2_n1867) );
  INV_X1 R2_U461 ( .A(R2_n1867), .ZN(R2_n1101) );
  AOI22_X1 R2_U460 ( .A1(n3335), .A2(R2_n2385), .B1(R2_n[688]), .B2(R2_n2382), 
        .ZN(R2_n1866) );
  INV_X1 R2_U459 ( .A(R2_n1866), .ZN(R2_n1102) );
  AOI22_X1 R2_U458 ( .A1(n3336), .A2(R2_n2384), .B1(R2_n[689]), .B2(R2_n2381), 
        .ZN(R2_n1865) );
  INV_X1 R2_U457 ( .A(R2_n1865), .ZN(R2_n1103) );
  AOI22_X1 R2_U456 ( .A1(n3337), .A2(R2_n2375), .B1(R2_n[690]), .B2(R2_n2379), 
        .ZN(R2_n1864) );
  INV_X1 R2_U455 ( .A(R2_n1864), .ZN(R2_n1104) );
  AOI22_X1 R2_U454 ( .A1(n3338), .A2(R2_n2383), .B1(R2_n[691]), .B2(R2_n2378), 
        .ZN(R2_n1863) );
  INV_X1 R2_U453 ( .A(R2_n1863), .ZN(R2_n1105) );
  AOI22_X1 R2_U452 ( .A1(n3339), .A2(R2_n2385), .B1(R2_n[692]), .B2(R2_n2377), 
        .ZN(R2_n1862) );
  INV_X1 R2_U451 ( .A(R2_n1862), .ZN(R2_n1106) );
  AOI22_X1 R2_U450 ( .A1(n3340), .A2(R2_n2375), .B1(R2_n[693]), .B2(R2_n2380), 
        .ZN(R2_n1861) );
  INV_X1 R2_U449 ( .A(R2_n1861), .ZN(R2_n1107) );
  AOI22_X1 R2_U448 ( .A1(n3341), .A2(R2_n2375), .B1(R2_n[694]), .B2(R2_n2379), 
        .ZN(R2_n1860) );
  INV_X1 R2_U447 ( .A(R2_n1860), .ZN(R2_n1108) );
  AOI22_X1 R2_U446 ( .A1(n3342), .A2(R2_n2375), .B1(R2_n[695]), .B2(R2_n2382), 
        .ZN(R2_n1859) );
  INV_X1 R2_U445 ( .A(R2_n1859), .ZN(R2_n1109) );
  AOI22_X1 R2_U444 ( .A1(n3343), .A2(R2_n2384), .B1(R2_n[696]), .B2(R2_n2381), 
        .ZN(R2_n1858) );
  INV_X1 R2_U443 ( .A(R2_n1858), .ZN(R2_n1110) );
  AOI22_X1 R2_U442 ( .A1(n3344), .A2(R2_n2375), .B1(R2_n[697]), .B2(R2_n2380), 
        .ZN(R2_n1857) );
  INV_X1 R2_U441 ( .A(R2_n1857), .ZN(R2_n1111) );
  AOI22_X1 R2_U440 ( .A1(n3345), .A2(R2_n2375), .B1(R2_n[698]), .B2(R2_n2380), 
        .ZN(R2_n1856) );
  INV_X1 R2_U439 ( .A(R2_n1856), .ZN(R2_n1112) );
  AOI22_X1 R2_U438 ( .A1(n3346), .A2(R2_n2376), .B1(R2_n[699]), .B2(R2_n2380), 
        .ZN(R2_n1855) );
  INV_X1 R2_U437 ( .A(R2_n1855), .ZN(R2_n1113) );
  AOI22_X1 R2_U436 ( .A1(n3347), .A2(R2_n2385), .B1(R2_n[700]), .B2(R2_n2380), 
        .ZN(R2_n1854) );
  INV_X1 R2_U435 ( .A(R2_n1854), .ZN(R2_n1114) );
  AOI22_X1 R2_U434 ( .A1(n3348), .A2(R2_n2383), .B1(R2_n[701]), .B2(R2_n2380), 
        .ZN(R2_n1853) );
  INV_X1 R2_U433 ( .A(R2_n1853), .ZN(R2_n1115) );
  AOI22_X1 R2_U432 ( .A1(n3349), .A2(R2_n2383), .B1(R2_n[702]), .B2(R2_n2380), 
        .ZN(R2_n1852) );
  INV_X1 R2_U431 ( .A(R2_n1852), .ZN(R2_n1116) );
  AOI22_X1 R2_U430 ( .A1(n3350), .A2(R2_n2384), .B1(R2_n[703]), .B2(R2_n2380), 
        .ZN(R2_n1851) );
  INV_X1 R2_U429 ( .A(R2_n1851), .ZN(R2_n1117) );
  AOI22_X1 R2_U428 ( .A1(n3351), .A2(R2_n2376), .B1(R2_n[704]), .B2(R2_n2380), 
        .ZN(R2_n1850) );
  INV_X1 R2_U427 ( .A(R2_n1850), .ZN(R2_n1118) );
  AOI22_X1 R2_U426 ( .A1(n3352), .A2(R2_n2384), .B1(R2_n[705]), .B2(R2_n2380), 
        .ZN(R2_n1849) );
  INV_X1 R2_U425 ( .A(R2_n1849), .ZN(R2_n1119) );
  AOI22_X1 R2_U424 ( .A1(n3353), .A2(R2_n2375), .B1(R2_n[706]), .B2(R2_n2379), 
        .ZN(R2_n1848) );
  INV_X1 R2_U423 ( .A(R2_n1848), .ZN(R2_n1120) );
  AOI22_X1 R2_U422 ( .A1(n3354), .A2(R2_n2375), .B1(R2_n[707]), .B2(R2_n2379), 
        .ZN(R2_n1847) );
  INV_X1 R2_U421 ( .A(R2_n1847), .ZN(R2_n1121) );
  AOI22_X1 R2_U420 ( .A1(n3355), .A2(R2_n1811), .B1(R2_n[708]), .B2(R2_n2379), 
        .ZN(R2_n1846) );
  INV_X1 R2_U419 ( .A(R2_n1846), .ZN(R2_n1122) );
  AOI22_X1 R2_U418 ( .A1(n3356), .A2(R2_n2383), .B1(R2_n[709]), .B2(R2_n2379), 
        .ZN(R2_n1845) );
  INV_X1 R2_U417 ( .A(R2_n1845), .ZN(R2_n1123) );
  AOI22_X1 R2_U416 ( .A1(n3357), .A2(R2_n2385), .B1(R2_n[710]), .B2(R2_n2379), 
        .ZN(R2_n1844) );
  INV_X1 R2_U415 ( .A(R2_n1844), .ZN(R2_n1124) );
  AOI22_X1 R2_U414 ( .A1(n3358), .A2(R2_n2383), .B1(R2_n[711]), .B2(R2_n2379), 
        .ZN(R2_n1843) );
  INV_X1 R2_U413 ( .A(R2_n1843), .ZN(R2_n1125) );
  AOI22_X1 R2_U412 ( .A1(n3359), .A2(R2_n2383), .B1(R2_n[712]), .B2(R2_n2379), 
        .ZN(R2_n1842) );
  INV_X1 R2_U411 ( .A(R2_n1842), .ZN(R2_n1126) );
  AOI22_X1 R2_U410 ( .A1(n3360), .A2(R2_n1811), .B1(R2_n[713]), .B2(R2_n2379), 
        .ZN(R2_n1841) );
  INV_X1 R2_U409 ( .A(R2_n1841), .ZN(R2_n1127) );
  AOI22_X1 R2_U408 ( .A1(n3361), .A2(R2_n2383), .B1(R2_n[714]), .B2(R2_n2379), 
        .ZN(R2_n1840) );
  INV_X1 R2_U407 ( .A(R2_n1840), .ZN(R2_n1128) );
  AOI22_X1 R2_U406 ( .A1(n3362), .A2(R2_n2385), .B1(R2_n[715]), .B2(R2_n2378), 
        .ZN(R2_n1839) );
  INV_X1 R2_U405 ( .A(R2_n1839), .ZN(R2_n1772) );
  AOI22_X1 R2_U404 ( .A1(n3363), .A2(R2_n2385), .B1(R2_n[716]), .B2(R2_n2378), 
        .ZN(R2_n1838) );
  INV_X1 R2_U403 ( .A(R2_n1838), .ZN(R2_n1773) );
  AOI22_X1 R2_U402 ( .A1(n3364), .A2(R2_n2385), .B1(R2_n[717]), .B2(R2_n2378), 
        .ZN(R2_n1837) );
  INV_X1 R2_U401 ( .A(R2_n1837), .ZN(R2_n1774) );
  AOI22_X1 R2_U400 ( .A1(n3365), .A2(R2_n2385), .B1(R2_n[718]), .B2(R2_n2378), 
        .ZN(R2_n1836) );
  INV_X1 R2_U399 ( .A(R2_n1836), .ZN(R2_n1775) );
  AOI22_X1 R2_U398 ( .A1(n3366), .A2(R2_n2383), .B1(R2_n[719]), .B2(R2_n2378), 
        .ZN(R2_n1835) );
  INV_X1 R2_U397 ( .A(R2_n1835), .ZN(R2_n1776) );
  AOI22_X1 R2_U396 ( .A1(n3367), .A2(R2_n2375), .B1(R2_n[720]), .B2(R2_n2378), 
        .ZN(R2_n1834) );
  INV_X1 R2_U395 ( .A(R2_n1834), .ZN(R2_n1777) );
  AOI22_X1 R2_U394 ( .A1(n3368), .A2(R2_n2383), .B1(R2_n[721]), .B2(R2_n2378), 
        .ZN(R2_n1833) );
  INV_X1 R2_U393 ( .A(R2_n1833), .ZN(R2_n1778) );
  AOI22_X1 R2_U392 ( .A1(n3369), .A2(R2_n2385), .B1(R2_n[722]), .B2(R2_n2378), 
        .ZN(R2_n1832) );
  INV_X1 R2_U391 ( .A(R2_n1832), .ZN(R2_n1779) );
  AOI22_X1 R2_U390 ( .A1(n3370), .A2(R2_n2384), .B1(R2_n[723]), .B2(R2_n2378), 
        .ZN(R2_n1831) );
  INV_X1 R2_U389 ( .A(R2_n1831), .ZN(R2_n1780) );
  AOI22_X1 R2_U388 ( .A1(n3371), .A2(R2_n2376), .B1(R2_n[724]), .B2(R2_n2382), 
        .ZN(R2_n1830) );
  INV_X1 R2_U387 ( .A(R2_n1830), .ZN(R2_n1781) );
  AOI22_X1 R2_U386 ( .A1(n3372), .A2(R2_n1811), .B1(R2_n[725]), .B2(R2_n2381), 
        .ZN(R2_n1829) );
  INV_X1 R2_U385 ( .A(R2_n1829), .ZN(R2_n1782) );
  AOI22_X1 R2_U384 ( .A1(n3373), .A2(R2_n2385), .B1(R2_n[726]), .B2(R2_n2382), 
        .ZN(R2_n1828) );
  INV_X1 R2_U383 ( .A(R2_n1828), .ZN(R2_n1783) );
  AOI22_X1 R2_U382 ( .A1(n3374), .A2(R2_n2375), .B1(R2_n[727]), .B2(R2_n2382), 
        .ZN(R2_n1827) );
  INV_X1 R2_U381 ( .A(R2_n1827), .ZN(R2_n1784) );
  AOI22_X1 R2_U380 ( .A1(n3375), .A2(R2_n2384), .B1(R2_n[728]), .B2(R2_n2382), 
        .ZN(R2_n1826) );
  INV_X1 R2_U379 ( .A(R2_n1826), .ZN(R2_n1785) );
  AOI22_X1 R2_U378 ( .A1(n3376), .A2(R2_n2384), .B1(R2_n[729]), .B2(R2_n2382), 
        .ZN(R2_n1825) );
  INV_X1 R2_U377 ( .A(R2_n1825), .ZN(R2_n1786) );
  AOI22_X1 R2_U376 ( .A1(n3377), .A2(R2_n2375), .B1(R2_n[730]), .B2(R2_n2382), 
        .ZN(R2_n1824) );
  INV_X1 R2_U375 ( .A(R2_n1824), .ZN(R2_n1787) );
  AOI22_X1 R2_U374 ( .A1(n3378), .A2(R2_n2375), .B1(R2_n[731]), .B2(R2_n2382), 
        .ZN(R2_n1823) );
  INV_X1 R2_U373 ( .A(R2_n1823), .ZN(R2_n1788) );
  AOI22_X1 R2_U372 ( .A1(n3379), .A2(R2_n2376), .B1(R2_n[732]), .B2(R2_n2382), 
        .ZN(R2_n1822) );
  INV_X1 R2_U371 ( .A(R2_n1822), .ZN(R2_n1789) );
  AOI22_X1 R2_U370 ( .A1(n3380), .A2(R2_n1811), .B1(R2_n[733]), .B2(R2_n2382), 
        .ZN(R2_n1821) );
  INV_X1 R2_U369 ( .A(R2_n1821), .ZN(R2_n1790) );
  AOI22_X1 R2_U368 ( .A1(n3381), .A2(R2_n2384), .B1(R2_n[734]), .B2(R2_n2382), 
        .ZN(R2_n1820) );
  INV_X1 R2_U367 ( .A(R2_n1820), .ZN(R2_n1791) );
  AOI22_X1 R2_U366 ( .A1(n3382), .A2(R2_n2376), .B1(R2_n[735]), .B2(R2_n2381), 
        .ZN(R2_n1819) );
  INV_X1 R2_U365 ( .A(R2_n1819), .ZN(R2_n1792) );
  AOI22_X1 R2_U364 ( .A1(n3383), .A2(R2_n2383), .B1(R2_n[736]), .B2(R2_n2381), 
        .ZN(R2_n1818) );
  INV_X1 R2_U363 ( .A(R2_n1818), .ZN(R2_n1793) );
  AOI22_X1 R2_U362 ( .A1(n3384), .A2(R2_n2376), .B1(R2_n[737]), .B2(R2_n2381), 
        .ZN(R2_n1817) );
  INV_X1 R2_U361 ( .A(R2_n1817), .ZN(R2_n1794) );
  AOI22_X1 R2_U360 ( .A1(n3385), .A2(R2_n2384), .B1(R2_n[738]), .B2(R2_n2381), 
        .ZN(R2_n1816) );
  INV_X1 R2_U359 ( .A(R2_n1816), .ZN(R2_n1795) );
  AOI22_X1 R2_U358 ( .A1(n3386), .A2(R2_n1811), .B1(R2_n[739]), .B2(R2_n2381), 
        .ZN(R2_n1815) );
  INV_X1 R2_U357 ( .A(R2_n1815), .ZN(R2_n1796) );
  AOI22_X1 R2_U356 ( .A1(n3387), .A2(R2_n2385), .B1(R2_n[740]), .B2(R2_n2381), 
        .ZN(R2_n1814) );
  INV_X1 R2_U355 ( .A(R2_n1814), .ZN(R2_n1797) );
  AOI22_X1 R2_U354 ( .A1(n3388), .A2(R2_n2375), .B1(R2_n[741]), .B2(R2_n2381), 
        .ZN(R2_n1813) );
  INV_X1 R2_U353 ( .A(R2_n1813), .ZN(R2_n1798) );
  AOI22_X1 R2_U352 ( .A1(n3389), .A2(R2_n2375), .B1(R2_n[742]), .B2(R2_n2381), 
        .ZN(R2_n1812) );
  INV_X1 R2_U351 ( .A(R2_n1812), .ZN(R2_n1799) );
  AOI22_X1 R2_U350 ( .A1(n3390), .A2(R2_n2375), .B1(R2_n[743]), .B2(R2_n2381), 
        .ZN(R2_n1810) );
  INV_X1 R2_U349 ( .A(R2_n1810), .ZN(R2_n1800) );
  AOI22_X1 R2_U348 ( .A1(R2_n2358), .A2(R2_n1258), .B1(R2_n2071), .B2(
        R2_U16_DATA1_0), .ZN(R2_n2198) );
  INV_X1 R2_U347 ( .A(R2_n2198), .ZN(R2_n131) );
  AOI22_X1 R2_U346 ( .A1(R2_n2358), .A2(R2_n1259), .B1(R2_n2364), .B2(
        R2_U16_DATA1_1), .ZN(R2_n2197) );
  INV_X1 R2_U345 ( .A(R2_n2197), .ZN(R2_n132) );
  AOI22_X1 R2_U344 ( .A1(R2_n2359), .A2(R2_n1260), .B1(R2_n2361), .B2(
        R2_U16_DATA1_2), .ZN(R2_n2196) );
  INV_X1 R2_U343 ( .A(R2_n2196), .ZN(R2_n133) );
  AOI22_X1 R2_U342 ( .A1(R2_n2358), .A2(R2_n1261), .B1(R2_n2361), .B2(
        R2_U16_DATA1_3), .ZN(R2_n2195) );
  INV_X1 R2_U341 ( .A(R2_n2195), .ZN(R2_n134) );
  AOI22_X1 R2_U340 ( .A1(R2_n2357), .A2(R2_n1262), .B1(R2_n2361), .B2(
        R2_U16_DATA1_4), .ZN(R2_n2194) );
  INV_X1 R2_U339 ( .A(R2_n2194), .ZN(R2_n135) );
  AOI22_X1 R2_U338 ( .A1(R2_n2358), .A2(R2_n1263), .B1(R2_n2071), .B2(
        R2_U16_DATA1_5), .ZN(R2_n2193) );
  INV_X1 R2_U337 ( .A(R2_n2193), .ZN(R2_n136) );
  AOI22_X1 R2_U336 ( .A1(R2_n2356), .A2(R2_n1264), .B1(R2_n2361), .B2(
        R2_U16_DATA1_6), .ZN(R2_n2192) );
  INV_X1 R2_U335 ( .A(R2_n2192), .ZN(R2_n137) );
  AOI22_X1 R2_U334 ( .A1(R2_n2355), .A2(R2_n1265), .B1(R2_n2364), .B2(
        R2_U16_DATA1_7), .ZN(R2_n2191) );
  INV_X1 R2_U333 ( .A(R2_n2191), .ZN(R2_n138) );
  INV_X1 R2_U331 ( .A(n3261), .ZN(R2_n1809) );
  OAI21_X1 R2_U330 ( .B1(n3261), .B2(R2_n1807), .A(R2_n2375), .ZN(R2_n2342) );
  NOR4_X1 R2_U329 ( .A1(R2_n1806), .A2(R2_r332_A_1_), .A3(R2_r332_A_2_), .A4(
        R2_r332_A_3_), .ZN(R2_n2333) );
  NOR4_X1 R2_U328 ( .A1(R2_n1805), .A2(R2_n1806), .A3(R2_r332_A_2_), .A4(
        R2_r332_A_3_), .ZN(R2_n2336) );
  AND2_X1 R2_U327 ( .A1(R2_n2331), .A2(R2_r332_A_3_), .ZN(R2_n2341) );
  AOI222_X1 R2_U326 ( .A1(R2_n260), .A2(R2_n2386), .B1(R2_U16_DATA2_35), .B2(
        R2_n2374), .C1(R2_U16_DATA1_35), .C2(R2_n2365), .ZN(R2_n2033) );
  INV_X1 R2_U325 ( .A(R2_n2033), .ZN(R2_n422) );
  AOI222_X1 R2_U324 ( .A1(R2_n261), .A2(R2_n2388), .B1(R2_U16_DATA2_36), .B2(
        R2_n2372), .C1(R2_U16_DATA1_36), .C2(R2_n1941), .ZN(R2_n2032) );
  INV_X1 R2_U323 ( .A(R2_n2032), .ZN(R2_n423) );
  AOI222_X1 R2_U322 ( .A1(R2_n262), .A2(R2_n2389), .B1(R2_U16_DATA2_37), .B2(
        R2_n2372), .C1(R2_U16_DATA1_37), .C2(R2_n1941), .ZN(R2_n2031) );
  INV_X1 R2_U321 ( .A(R2_n2031), .ZN(R2_n424) );
  AOI222_X1 R2_U320 ( .A1(R2_n263), .A2(R2_n2386), .B1(R2_U16_DATA2_38), .B2(
        R2_n2372), .C1(R2_U16_DATA1_38), .C2(R2_n1941), .ZN(R2_n2030) );
  INV_X1 R2_U319 ( .A(R2_n2030), .ZN(R2_n425) );
  AOI222_X1 R2_U318 ( .A1(R2_n264), .A2(R2_n2390), .B1(R2_U16_DATA2_39), .B2(
        R2_n2372), .C1(R2_U16_DATA1_39), .C2(R2_n1941), .ZN(R2_n2029) );
  INV_X1 R2_U317 ( .A(R2_n2029), .ZN(R2_n426) );
  AOI222_X1 R2_U316 ( .A1(R2_n265), .A2(R2_n2387), .B1(R2_U16_DATA2_40), .B2(
        R2_n2372), .C1(R2_U16_DATA1_40), .C2(R2_n1941), .ZN(R2_n2028) );
  INV_X1 R2_U315 ( .A(R2_n2028), .ZN(R2_n427) );
  AOI222_X1 R2_U314 ( .A1(R2_n266), .A2(R2_n2388), .B1(R2_U16_DATA2_41), .B2(
        R2_n2372), .C1(R2_U16_DATA1_41), .C2(R2_n1941), .ZN(R2_n2027) );
  INV_X1 R2_U313 ( .A(R2_n2027), .ZN(R2_n428) );
  AOI222_X1 R2_U312 ( .A1(R2_n267), .A2(R2_n2389), .B1(R2_U16_DATA2_42), .B2(
        R2_n2372), .C1(R2_U16_DATA1_42), .C2(R2_n1941), .ZN(R2_n2026) );
  INV_X1 R2_U311 ( .A(R2_n2026), .ZN(R2_n429) );
  AOI222_X1 R2_U310 ( .A1(R2_n268), .A2(R2_n2386), .B1(R2_U16_DATA2_43), .B2(
        R2_n2372), .C1(R2_U16_DATA1_43), .C2(R2_n2365), .ZN(R2_n2025) );
  INV_X1 R2_U309 ( .A(R2_n2025), .ZN(R2_n430) );
  AOI222_X1 R2_U308 ( .A1(R2_n269), .A2(R2_n2390), .B1(R2_U16_DATA2_44), .B2(
        R2_n2372), .C1(R2_U16_DATA1_44), .C2(R2_n2369), .ZN(R2_n2024) );
  INV_X1 R2_U307 ( .A(R2_n2024), .ZN(R2_n431) );
  AOI222_X1 R2_U306 ( .A1(R2_n270), .A2(R2_n2387), .B1(R2_U16_DATA2_45), .B2(
        R2_n2372), .C1(R2_U16_DATA1_45), .C2(R2_n2365), .ZN(R2_n2023) );
  INV_X1 R2_U305 ( .A(R2_n2023), .ZN(R2_n432) );
  AOI222_X1 R2_U304 ( .A1(R2_n271), .A2(R2_n2388), .B1(R2_U16_DATA2_46), .B2(
        R2_n2372), .C1(R2_U16_DATA1_46), .C2(R2_n2365), .ZN(R2_n2022) );
  INV_X1 R2_U303 ( .A(R2_n2022), .ZN(R2_n433) );
  AOI222_X1 R2_U302 ( .A1(R2_n272), .A2(R2_n2386), .B1(R2_U16_DATA2_47), .B2(
        R2_n2372), .C1(R2_U16_DATA1_47), .C2(R2_n2365), .ZN(R2_n2021) );
  INV_X1 R2_U301 ( .A(R2_n2021), .ZN(R2_n434) );
  AOI222_X1 R2_U300 ( .A1(R2_n273), .A2(R2_n2387), .B1(R2_U16_DATA2_48), .B2(
        R2_n2373), .C1(R2_U16_DATA1_48), .C2(R2_n1941), .ZN(R2_n2020) );
  INV_X1 R2_U299 ( .A(R2_n2020), .ZN(R2_n435) );
  AOI222_X1 R2_U298 ( .A1(R2_n274), .A2(R2_n2388), .B1(R2_U16_DATA2_49), .B2(
        R2_n2373), .C1(R2_U16_DATA1_49), .C2(R2_n1941), .ZN(R2_n2019) );
  INV_X1 R2_U297 ( .A(R2_n2019), .ZN(R2_n436) );
  AOI222_X1 R2_U296 ( .A1(R2_n275), .A2(R2_n2389), .B1(R2_U16_DATA2_50), .B2(
        R2_n2373), .C1(R2_U16_DATA1_50), .C2(R2_n1941), .ZN(R2_n2018) );
  INV_X1 R2_U295 ( .A(R2_n2018), .ZN(R2_n437) );
  AOI222_X1 R2_U294 ( .A1(R2_n276), .A2(R2_n2386), .B1(R2_U16_DATA2_51), .B2(
        R2_n2373), .C1(R2_U16_DATA1_51), .C2(R2_n1941), .ZN(R2_n2017) );
  INV_X1 R2_U293 ( .A(R2_n2017), .ZN(R2_n438) );
  AOI222_X1 R2_U292 ( .A1(R2_n277), .A2(R2_n2387), .B1(R2_U16_DATA2_52), .B2(
        R2_n2373), .C1(R2_U16_DATA1_52), .C2(R2_n1941), .ZN(R2_n2016) );
  INV_X1 R2_U291 ( .A(R2_n2016), .ZN(R2_n439) );
  AOI222_X1 R2_U290 ( .A1(R2_n278), .A2(R2_n2388), .B1(R2_U16_DATA2_53), .B2(
        R2_n2373), .C1(R2_U16_DATA1_53), .C2(R2_n1941), .ZN(R2_n2015) );
  INV_X1 R2_U289 ( .A(R2_n2015), .ZN(R2_n440) );
  AOI222_X1 R2_U288 ( .A1(R2_n279), .A2(R2_n2389), .B1(R2_U16_DATA2_54), .B2(
        R2_n2373), .C1(R2_U16_DATA1_54), .C2(R2_n1941), .ZN(R2_n2014) );
  INV_X1 R2_U287 ( .A(R2_n2014), .ZN(R2_n441) );
  AOI222_X1 R2_U286 ( .A1(R2_n280), .A2(R2_n2386), .B1(R2_U16_DATA2_55), .B2(
        R2_n2373), .C1(R2_U16_DATA1_55), .C2(R2_n1941), .ZN(R2_n2013) );
  INV_X1 R2_U285 ( .A(R2_n2013), .ZN(R2_n442) );
  AOI222_X1 R2_U284 ( .A1(R2_n281), .A2(R2_n2387), .B1(R2_U16_DATA2_56), .B2(
        R2_n2373), .C1(R2_U16_DATA1_56), .C2(R2_n2365), .ZN(R2_n2012) );
  INV_X1 R2_U283 ( .A(R2_n2012), .ZN(R2_n443) );
  AOI222_X1 R2_U282 ( .A1(R2_n282), .A2(R2_n2388), .B1(R2_U16_DATA2_57), .B2(
        R2_n2373), .C1(R2_U16_DATA1_57), .C2(R2_n2368), .ZN(R2_n2011) );
  INV_X1 R2_U281 ( .A(R2_n2011), .ZN(R2_n444) );
  AOI222_X1 R2_U280 ( .A1(R2_n283), .A2(R2_n2389), .B1(R2_U16_DATA2_58), .B2(
        R2_n2373), .C1(R2_U16_DATA1_58), .C2(R2_n2365), .ZN(R2_n2010) );
  INV_X1 R2_U279 ( .A(R2_n2010), .ZN(R2_n445) );
  AOI222_X1 R2_U278 ( .A1(R2_n284), .A2(R2_n2386), .B1(R2_U16_DATA2_59), .B2(
        R2_n2373), .C1(R2_U16_DATA1_59), .C2(R2_n2365), .ZN(R2_n2009) );
  INV_X1 R2_U277 ( .A(R2_n2009), .ZN(R2_n446) );
  AOI222_X1 R2_U276 ( .A1(R2_n285), .A2(R2_n2390), .B1(R2_U16_DATA2_60), .B2(
        R2_n2374), .C1(R2_U16_DATA1_60), .C2(R2_n2365), .ZN(R2_n2008) );
  INV_X1 R2_U275 ( .A(R2_n2008), .ZN(R2_n447) );
  AOI222_X1 R2_U274 ( .A1(R2_n286), .A2(R2_n2390), .B1(R2_U16_DATA2_61), .B2(
        R2_n2374), .C1(R2_U16_DATA1_61), .C2(R2_n2367), .ZN(R2_n2007) );
  INV_X1 R2_U273 ( .A(R2_n2007), .ZN(R2_n448) );
  AOI222_X1 R2_U272 ( .A1(R2_n287), .A2(R2_n2390), .B1(R2_U16_DATA2_62), .B2(
        R2_n2374), .C1(R2_U16_DATA1_62), .C2(R2_n2365), .ZN(R2_n2006) );
  INV_X1 R2_U271 ( .A(R2_n2006), .ZN(R2_n449) );
  AOI222_X1 R2_U270 ( .A1(R2_n288), .A2(R2_n2390), .B1(R2_U16_DATA2_63), .B2(
        R2_n2374), .C1(R2_U16_DATA1_63), .C2(R2_n2365), .ZN(R2_n2005) );
  INV_X1 R2_U269 ( .A(R2_n2005), .ZN(R2_n450) );
  AOI222_X1 R2_U268 ( .A1(R2_n289), .A2(R2_n2390), .B1(R2_U16_DATA2_64), .B2(
        R2_n2374), .C1(R2_U16_DATA1_64), .C2(R2_n2368), .ZN(R2_n2004) );
  INV_X1 R2_U267 ( .A(R2_n2004), .ZN(R2_n451) );
  AOI222_X1 R2_U266 ( .A1(R2_n290), .A2(R2_n2390), .B1(R2_U16_DATA2_65), .B2(
        R2_n2374), .C1(R2_U16_DATA1_65), .C2(R2_n1941), .ZN(R2_n2003) );
  INV_X1 R2_U265 ( .A(R2_n2003), .ZN(R2_n452) );
  AOI222_X1 R2_U264 ( .A1(R2_n291), .A2(R2_n2390), .B1(R2_U16_DATA2_66), .B2(
        R2_n2374), .C1(R2_U16_DATA1_66), .C2(R2_n1941), .ZN(R2_n2002) );
  INV_X1 R2_U263 ( .A(R2_n2002), .ZN(R2_n453) );
  AOI222_X1 R2_U262 ( .A1(R2_n292), .A2(R2_n2386), .B1(R2_U16_DATA2_67), .B2(
        R2_n2374), .C1(R2_U16_DATA1_67), .C2(R2_n1941), .ZN(R2_n2001) );
  INV_X1 R2_U261 ( .A(R2_n2001), .ZN(R2_n454) );
  AOI222_X1 R2_U260 ( .A1(R2_n293), .A2(R2_n2386), .B1(R2_U16_DATA2_68), .B2(
        R2_n2374), .C1(R2_U16_DATA1_68), .C2(R2_n2365), .ZN(R2_n2000) );
  INV_X1 R2_U259 ( .A(R2_n2000), .ZN(R2_n455) );
  AOI222_X1 R2_U258 ( .A1(R2_n294), .A2(R2_n2386), .B1(R2_U16_DATA2_69), .B2(
        R2_n2374), .C1(R2_U16_DATA1_69), .C2(R2_n2365), .ZN(R2_n1999) );
  INV_X1 R2_U257 ( .A(R2_n1999), .ZN(R2_n456) );
  AOI222_X1 R2_U256 ( .A1(R2_n295), .A2(R2_n2386), .B1(R2_U16_DATA2_70), .B2(
        R2_n2374), .C1(R2_U16_DATA1_70), .C2(R2_n2369), .ZN(R2_n1998) );
  INV_X1 R2_U255 ( .A(R2_n1998), .ZN(R2_n457) );
  AOI222_X1 R2_U254 ( .A1(R2_n320), .A2(R2_n2389), .B1(R2_U16_DATA2_95), .B2(
        R2_n1940), .C1(R2_U16_DATA1_95), .C2(R2_n2367), .ZN(R2_n1973) );
  INV_X1 R2_U253 ( .A(R2_n1973), .ZN(R2_n611) );
  AOI222_X1 R2_U252 ( .A1(R2_n321), .A2(R2_n2389), .B1(R2_U16_DATA2_96), .B2(
        R2_n1940), .C1(R2_U16_DATA1_96), .C2(R2_n1941), .ZN(R2_n1972) );
  INV_X1 R2_U251 ( .A(R2_n1972), .ZN(R2_n612) );
  AOI222_X1 R2_U250 ( .A1(R2_n322), .A2(R2_n2389), .B1(R2_U16_DATA2_97), .B2(
        R2_n1940), .C1(R2_U16_DATA1_97), .C2(R2_n1941), .ZN(R2_n1971) );
  INV_X1 R2_U249 ( .A(R2_n1971), .ZN(R2_n613) );
  AOI222_X1 R2_U248 ( .A1(R2_n323), .A2(R2_n2389), .B1(R2_U16_DATA2_98), .B2(
        R2_n1940), .C1(R2_U16_DATA1_98), .C2(R2_n1941), .ZN(R2_n1970) );
  INV_X1 R2_U247 ( .A(R2_n1970), .ZN(R2_n614) );
  AOI222_X1 R2_U246 ( .A1(R2_n324), .A2(R2_n2389), .B1(R2_U16_DATA2_99), .B2(
        R2_n2370), .C1(R2_U16_DATA1_99), .C2(R2_n1941), .ZN(R2_n1969) );
  INV_X1 R2_U245 ( .A(R2_n1969), .ZN(R2_n1001) );
  AOI222_X1 R2_U244 ( .A1(R2_n325), .A2(R2_n2389), .B1(R2_U16_DATA2_100), .B2(
        R2_n2370), .C1(R2_U16_DATA1_100), .C2(R2_n2368), .ZN(R2_n1968) );
  INV_X1 R2_U243 ( .A(R2_n1968), .ZN(R2_n1002) );
  AOI222_X1 R2_U242 ( .A1(R2_n326), .A2(R2_n2389), .B1(R2_U16_DATA2_101), .B2(
        R2_n2370), .C1(R2_U16_DATA1_101), .C2(R2_n2365), .ZN(R2_n1967) );
  INV_X1 R2_U241 ( .A(R2_n1967), .ZN(R2_n1003) );
  AOI222_X1 R2_U240 ( .A1(R2_n327), .A2(R2_n2389), .B1(R2_U16_DATA2_102), .B2(
        R2_n2370), .C1(R2_U16_DATA1_102), .C2(R2_n2369), .ZN(R2_n1966) );
  INV_X1 R2_U239 ( .A(R2_n1966), .ZN(R2_n1004) );
  AOI222_X1 R2_U238 ( .A1(R2_n328), .A2(R2_n2389), .B1(R2_U16_DATA2_103), .B2(
        R2_n2371), .C1(R2_U16_DATA1_103), .C2(R2_n2366), .ZN(R2_n1965) );
  INV_X1 R2_U237 ( .A(R2_n1965), .ZN(R2_n1005) );
  AOI222_X1 R2_U236 ( .A1(R2_n329), .A2(R2_n2389), .B1(R2_U16_DATA2_104), .B2(
        R2_n2370), .C1(R2_U16_DATA1_104), .C2(R2_n2369), .ZN(R2_n1964) );
  INV_X1 R2_U235 ( .A(R2_n1964), .ZN(R2_n1006) );
  AOI222_X1 R2_U234 ( .A1(R2_n330), .A2(R2_n2389), .B1(R2_U16_DATA2_105), .B2(
        R2_n2370), .C1(R2_U16_DATA1_105), .C2(R2_n2369), .ZN(R2_n1963) );
  INV_X1 R2_U233 ( .A(R2_n1963), .ZN(R2_n1007) );
  AOI222_X1 R2_U232 ( .A1(R2_n331), .A2(R2_n2389), .B1(R2_U16_DATA2_106), .B2(
        R2_n2371), .C1(R2_U16_DATA1_106), .C2(R2_n2369), .ZN(R2_n1962) );
  INV_X1 R2_U231 ( .A(R2_n1962), .ZN(R2_n1008) );
  AOI222_X1 R2_U230 ( .A1(R2_n332), .A2(R2_n2387), .B1(R2_U16_DATA2_107), .B2(
        R2_n2371), .C1(R2_U16_DATA1_107), .C2(R2_n2369), .ZN(R2_n1961) );
  INV_X1 R2_U229 ( .A(R2_n1961), .ZN(R2_n1009) );
  AOI222_X1 R2_U228 ( .A1(R2_n333), .A2(R2_n2386), .B1(R2_U16_DATA2_108), .B2(
        R2_n2370), .C1(R2_U16_DATA1_108), .C2(R2_n2368), .ZN(R2_n1960) );
  INV_X1 R2_U227 ( .A(R2_n1960), .ZN(R2_n1010) );
  AOI222_X1 R2_U226 ( .A1(R2_n334), .A2(R2_n2389), .B1(R2_U16_DATA2_109), .B2(
        R2_n2370), .C1(R2_U16_DATA1_109), .C2(R2_n2368), .ZN(R2_n1959) );
  INV_X1 R2_U225 ( .A(R2_n1959), .ZN(R2_n1011) );
  AOI222_X1 R2_U224 ( .A1(R2_n335), .A2(R2_n2386), .B1(R2_U16_DATA2_110), .B2(
        R2_n2371), .C1(R2_U16_DATA1_110), .C2(R2_n2368), .ZN(R2_n1958) );
  INV_X1 R2_U223 ( .A(R2_n1958), .ZN(R2_n1012) );
  AOI222_X1 R2_U222 ( .A1(R2_n336), .A2(R2_n2387), .B1(R2_U16_DATA2_111), .B2(
        R2_n2371), .C1(R2_U16_DATA1_111), .C2(R2_n2368), .ZN(R2_n1957) );
  INV_X1 R2_U221 ( .A(R2_n1957), .ZN(R2_n1013) );
  AOI222_X1 R2_U220 ( .A1(R2_n337), .A2(R2_n2386), .B1(R2_U16_DATA2_112), .B2(
        R2_n2370), .C1(R2_U16_DATA1_112), .C2(R2_n2368), .ZN(R2_n1956) );
  INV_X1 R2_U219 ( .A(R2_n1956), .ZN(R2_n1014) );
  AOI222_X1 R2_U218 ( .A1(R2_n338), .A2(R2_n2388), .B1(R2_U16_DATA2_113), .B2(
        R2_n2370), .C1(R2_U16_DATA1_113), .C2(R2_n2368), .ZN(R2_n1955) );
  INV_X1 R2_U217 ( .A(R2_n1955), .ZN(R2_n1015) );
  AOI222_X1 R2_U216 ( .A1(R2_n339), .A2(R2_n2386), .B1(R2_U16_DATA2_114), .B2(
        R2_n2371), .C1(R2_U16_DATA1_114), .C2(R2_n2368), .ZN(R2_n1954) );
  INV_X1 R2_U215 ( .A(R2_n1954), .ZN(R2_n1016) );
  AOI222_X1 R2_U214 ( .A1(R2_n340), .A2(R2_n2389), .B1(R2_U16_DATA2_115), .B2(
        R2_n2371), .C1(R2_U16_DATA1_115), .C2(R2_n2368), .ZN(R2_n1953) );
  INV_X1 R2_U213 ( .A(R2_n1953), .ZN(R2_n1017) );
  AOI222_X1 R2_U212 ( .A1(R2_n341), .A2(R2_n2386), .B1(R2_U16_DATA2_116), .B2(
        R2_n2370), .C1(R2_U16_DATA1_116), .C2(R2_n2368), .ZN(R2_n1952) );
  INV_X1 R2_U211 ( .A(R2_n1952), .ZN(R2_n1018) );
  AOI222_X1 R2_U210 ( .A1(R2_n342), .A2(R2_n2387), .B1(R2_U16_DATA2_117), .B2(
        R2_n2370), .C1(R2_U16_DATA1_117), .C2(R2_n2368), .ZN(R2_n1951) );
  INV_X1 R2_U209 ( .A(R2_n1951), .ZN(R2_n1019) );
  AOI222_X1 R2_U208 ( .A1(R2_n343), .A2(R2_n2388), .B1(R2_U16_DATA2_118), .B2(
        R2_n2370), .C1(R2_U16_DATA1_118), .C2(R2_n2368), .ZN(R2_n1950) );
  INV_X1 R2_U207 ( .A(R2_n1950), .ZN(R2_n1020) );
  AOI222_X1 R2_U206 ( .A1(R2_n344), .A2(R2_n2390), .B1(R2_U16_DATA2_119), .B2(
        R2_n2373), .C1(R2_U16_DATA1_119), .C2(R2_n2368), .ZN(R2_n1949) );
  INV_X1 R2_U205 ( .A(R2_n1949), .ZN(R2_n1021) );
  AOI222_X1 R2_U204 ( .A1(R2_n345), .A2(R2_n2390), .B1(R2_U16_DATA2_120), .B2(
        R2_n2373), .C1(R2_U16_DATA1_120), .C2(R2_n2369), .ZN(R2_n1948) );
  INV_X1 R2_U203 ( .A(R2_n1948), .ZN(R2_n1022) );
  AOI222_X1 R2_U202 ( .A1(R2_n346), .A2(R2_n2390), .B1(R2_U16_DATA2_121), .B2(
        R2_n2373), .C1(R2_U16_DATA1_121), .C2(R2_n2369), .ZN(R2_n1947) );
  INV_X1 R2_U201 ( .A(R2_n1947), .ZN(R2_n1023) );
  AOI222_X1 R2_U200 ( .A1(R2_n347), .A2(R2_n2390), .B1(R2_U16_DATA2_122), .B2(
        R2_n2373), .C1(R2_U16_DATA1_122), .C2(R2_n2369), .ZN(R2_n1946) );
  INV_X1 R2_U199 ( .A(R2_n1946), .ZN(R2_n1024) );
  AOI222_X1 R2_U198 ( .A1(R2_n348), .A2(R2_n2390), .B1(R2_U16_DATA2_123), .B2(
        R2_n2373), .C1(R2_U16_DATA1_123), .C2(R2_n2369), .ZN(R2_n1945) );
  INV_X1 R2_U197 ( .A(R2_n1945), .ZN(R2_n1025) );
  AOI222_X1 R2_U196 ( .A1(R2_n349), .A2(R2_n2390), .B1(R2_U16_DATA2_124), .B2(
        R2_n2373), .C1(R2_U16_DATA1_124), .C2(R2_n2369), .ZN(R2_n1944) );
  INV_X1 R2_U195 ( .A(R2_n1944), .ZN(R2_n1026) );
  AOI222_X1 R2_U194 ( .A1(R2_n350), .A2(R2_n2390), .B1(R2_U16_DATA2_125), .B2(
        R2_n2373), .C1(R2_U16_DATA1_125), .C2(R2_n2369), .ZN(R2_n1943) );
  INV_X1 R2_U193 ( .A(R2_n1943), .ZN(R2_n1027) );
  AOI222_X1 R2_U192 ( .A1(R2_n351), .A2(R2_n2390), .B1(R2_U16_DATA2_126), .B2(
        R2_n2370), .C1(R2_U16_DATA1_126), .C2(R2_n2369), .ZN(R2_n1942) );
  INV_X1 R2_U191 ( .A(R2_n1942), .ZN(R2_n1028) );
  AOI222_X1 R2_U190 ( .A1(R2_n352), .A2(R2_n2390), .B1(R2_U16_DATA2_127), .B2(
        R2_n2370), .C1(R2_U16_DATA1_127), .C2(R2_n2369), .ZN(R2_n1939) );
  INV_X1 R2_U189 ( .A(R2_n1939), .ZN(R2_n1029) );
  AOI222_X1 R2_U188 ( .A1(R2_n225), .A2(R2_n1802), .B1(R2_U16_DATA2_0), .B2(
        R2_n2371), .C1(R2_U16_DATA1_0), .C2(R2_n2365), .ZN(R2_n2068) );
  INV_X1 R2_U187 ( .A(R2_n2068), .ZN(R2_n387) );
  AOI222_X1 R2_U186 ( .A1(R2_n226), .A2(R2_n1802), .B1(R2_U16_DATA2_1), .B2(
        R2_n2371), .C1(R2_U16_DATA1_1), .C2(R2_n2365), .ZN(R2_n2067) );
  INV_X1 R2_U185 ( .A(R2_n2067), .ZN(R2_n388) );
  AOI222_X1 R2_U184 ( .A1(R2_n227), .A2(R2_n1802), .B1(R2_U16_DATA2_2), .B2(
        R2_n2370), .C1(R2_U16_DATA1_2), .C2(R2_n2368), .ZN(R2_n2066) );
  INV_X1 R2_U183 ( .A(R2_n2066), .ZN(R2_n389) );
  AOI222_X1 R2_U182 ( .A1(R2_n228), .A2(R2_n1802), .B1(R2_U16_DATA2_3), .B2(
        R2_n2370), .C1(R2_U16_DATA1_3), .C2(R2_n2366), .ZN(R2_n2065) );
  INV_X1 R2_U181 ( .A(R2_n2065), .ZN(R2_n390) );
  AOI222_X1 R2_U180 ( .A1(R2_n229), .A2(R2_n1802), .B1(R2_U16_DATA2_4), .B2(
        R2_n2371), .C1(R2_U16_DATA1_4), .C2(R2_n2365), .ZN(R2_n2064) );
  INV_X1 R2_U179 ( .A(R2_n2064), .ZN(R2_n391) );
  AOI222_X1 R2_U178 ( .A1(R2_n230), .A2(R2_n1802), .B1(R2_U16_DATA2_5), .B2(
        R2_n2370), .C1(R2_U16_DATA1_5), .C2(R2_n2365), .ZN(R2_n2063) );
  INV_X1 R2_U177 ( .A(R2_n2063), .ZN(R2_n392) );
  AOI222_X1 R2_U176 ( .A1(R2_n231), .A2(R2_n1802), .B1(R2_U16_DATA2_6), .B2(
        R2_n2371), .C1(R2_U16_DATA1_6), .C2(R2_n2365), .ZN(R2_n2062) );
  INV_X1 R2_U175 ( .A(R2_n2062), .ZN(R2_n393) );
  AOI222_X1 R2_U174 ( .A1(R2_n232), .A2(R2_n1802), .B1(R2_U16_DATA2_7), .B2(
        R2_n2371), .C1(R2_U16_DATA1_7), .C2(R2_n1941), .ZN(R2_n2061) );
  INV_X1 R2_U173 ( .A(R2_n2061), .ZN(R2_n394) );
  AOI222_X1 R2_U172 ( .A1(R2_n233), .A2(R2_n1802), .B1(R2_U16_DATA2_8), .B2(
        R2_n2370), .C1(R2_U16_DATA1_8), .C2(R2_n2369), .ZN(R2_n2060) );
  INV_X1 R2_U171 ( .A(R2_n2060), .ZN(R2_n395) );
  AOI222_X1 R2_U170 ( .A1(R2_n234), .A2(R2_n1802), .B1(R2_U16_DATA2_9), .B2(
        R2_n2371), .C1(R2_U16_DATA1_9), .C2(R2_n2366), .ZN(R2_n2059) );
  INV_X1 R2_U169 ( .A(R2_n2059), .ZN(R2_n396) );
  AOI222_X1 R2_U168 ( .A1(R2_n235), .A2(R2_n1802), .B1(R2_U16_DATA2_10), .B2(
        R2_n2371), .C1(R2_U16_DATA1_10), .C2(R2_n2365), .ZN(R2_n2058) );
  INV_X1 R2_U167 ( .A(R2_n2058), .ZN(R2_n397) );
  AOI222_X1 R2_U166 ( .A1(R2_n236), .A2(R2_n2386), .B1(R2_U16_DATA2_11), .B2(
        R2_n2370), .C1(R2_U16_DATA1_11), .C2(R2_n2365), .ZN(R2_n2057) );
  INV_X1 R2_U165 ( .A(R2_n2057), .ZN(R2_n398) );
  AOI222_X1 R2_U164 ( .A1(R2_n237), .A2(R2_n2387), .B1(R2_U16_DATA2_12), .B2(
        R2_n2372), .C1(R2_U16_DATA1_12), .C2(R2_n2367), .ZN(R2_n2056) );
  INV_X1 R2_U163 ( .A(R2_n2056), .ZN(R2_n399) );
  AOI222_X1 R2_U162 ( .A1(R2_n238), .A2(R2_n2390), .B1(R2_U16_DATA2_13), .B2(
        R2_n2374), .C1(R2_U16_DATA1_13), .C2(R2_n2367), .ZN(R2_n2055) );
  INV_X1 R2_U161 ( .A(R2_n2055), .ZN(R2_n400) );
  AOI222_X1 R2_U160 ( .A1(R2_n239), .A2(R2_n2389), .B1(R2_U16_DATA2_14), .B2(
        R2_n2372), .C1(R2_U16_DATA1_14), .C2(R2_n2365), .ZN(R2_n2054) );
  INV_X1 R2_U159 ( .A(R2_n2054), .ZN(R2_n401) );
  AOI222_X1 R2_U158 ( .A1(R2_n240), .A2(R2_n2388), .B1(R2_U16_DATA2_15), .B2(
        R2_n2372), .C1(R2_U16_DATA1_15), .C2(R2_n2365), .ZN(R2_n2053) );
  INV_X1 R2_U157 ( .A(R2_n2053), .ZN(R2_n402) );
  AOI222_X1 R2_U156 ( .A1(R2_n241), .A2(R2_n2389), .B1(R2_U16_DATA2_16), .B2(
        R2_n2374), .C1(R2_U16_DATA1_16), .C2(R2_n2365), .ZN(R2_n2052) );
  INV_X1 R2_U155 ( .A(R2_n2052), .ZN(R2_n403) );
  AOI222_X1 R2_U154 ( .A1(R2_n242), .A2(R2_n2388), .B1(R2_U16_DATA2_17), .B2(
        R2_n2374), .C1(R2_U16_DATA1_17), .C2(R2_n2365), .ZN(R2_n2051) );
  INV_X1 R2_U153 ( .A(R2_n2051), .ZN(R2_n404) );
  AOI222_X1 R2_U152 ( .A1(R2_n243), .A2(R2_n2387), .B1(R2_U16_DATA2_18), .B2(
        R2_n2372), .C1(R2_U16_DATA1_18), .C2(R2_n2368), .ZN(R2_n2050) );
  INV_X1 R2_U151 ( .A(R2_n2050), .ZN(R2_n405) );
  AOI222_X1 R2_U150 ( .A1(R2_n244), .A2(R2_n2386), .B1(R2_U16_DATA2_19), .B2(
        R2_n2374), .C1(R2_U16_DATA1_19), .C2(R2_n2368), .ZN(R2_n2049) );
  INV_X1 R2_U149 ( .A(R2_n2049), .ZN(R2_n406) );
  AOI222_X1 R2_U148 ( .A1(R2_n245), .A2(R2_n2390), .B1(R2_U16_DATA2_20), .B2(
        R2_n2372), .C1(R2_U16_DATA1_20), .C2(R2_n2365), .ZN(R2_n2048) );
  INV_X1 R2_U147 ( .A(R2_n2048), .ZN(R2_n407) );
  AOI222_X1 R2_U146 ( .A1(R2_n246), .A2(R2_n2386), .B1(R2_U16_DATA2_21), .B2(
        R2_n2372), .C1(R2_U16_DATA1_21), .C2(R2_n2365), .ZN(R2_n2047) );
  INV_X1 R2_U145 ( .A(R2_n2047), .ZN(R2_n408) );
  AOI222_X1 R2_U144 ( .A1(R2_n247), .A2(R2_n2386), .B1(R2_U16_DATA2_22), .B2(
        R2_n2371), .C1(R2_U16_DATA1_22), .C2(R2_n2365), .ZN(R2_n2046) );
  INV_X1 R2_U143 ( .A(R2_n2046), .ZN(R2_n409) );
  AOI222_X1 R2_U142 ( .A1(R2_n248), .A2(R2_n2390), .B1(R2_U16_DATA2_23), .B2(
        R2_n2371), .C1(R2_U16_DATA1_23), .C2(R2_n2365), .ZN(R2_n2045) );
  INV_X1 R2_U141 ( .A(R2_n2045), .ZN(R2_n410) );
  AOI222_X1 R2_U140 ( .A1(R2_n249), .A2(R2_n2389), .B1(R2_U16_DATA2_24), .B2(
        R2_n2372), .C1(R2_U16_DATA1_24), .C2(R2_n2365), .ZN(R2_n2044) );
  INV_X1 R2_U139 ( .A(R2_n2044), .ZN(R2_n411) );
  AOI222_X1 R2_U138 ( .A1(R2_n250), .A2(R2_n2390), .B1(R2_U16_DATA2_25), .B2(
        R2_n2374), .C1(R2_U16_DATA1_25), .C2(R2_n2365), .ZN(R2_n2043) );
  INV_X1 R2_U137 ( .A(R2_n2043), .ZN(R2_n412) );
  AOI222_X1 R2_U136 ( .A1(R2_n251), .A2(R2_n2388), .B1(R2_U16_DATA2_26), .B2(
        R2_n2372), .C1(R2_U16_DATA1_26), .C2(R2_n2365), .ZN(R2_n2042) );
  INV_X1 R2_U135 ( .A(R2_n2042), .ZN(R2_n413) );
  AOI222_X1 R2_U134 ( .A1(R2_n252), .A2(R2_n2387), .B1(R2_U16_DATA2_27), .B2(
        R2_n2374), .C1(R2_U16_DATA1_27), .C2(R2_n2365), .ZN(R2_n2041) );
  INV_X1 R2_U133 ( .A(R2_n2041), .ZN(R2_n414) );
  AOI222_X1 R2_U132 ( .A1(R2_n253), .A2(R2_n2387), .B1(R2_U16_DATA2_28), .B2(
        R2_n2372), .C1(R2_U16_DATA1_28), .C2(R2_n2365), .ZN(R2_n2040) );
  INV_X1 R2_U131 ( .A(R2_n2040), .ZN(R2_n415) );
  AOI222_X1 R2_U130 ( .A1(R2_n254), .A2(R2_n2389), .B1(R2_U16_DATA2_29), .B2(
        R2_n2374), .C1(R2_U16_DATA1_29), .C2(R2_n2365), .ZN(R2_n2039) );
  INV_X1 R2_U129 ( .A(R2_n2039), .ZN(R2_n416) );
  AOI222_X1 R2_U128 ( .A1(R2_n255), .A2(R2_n2388), .B1(R2_U16_DATA2_30), .B2(
        R2_n2374), .C1(R2_U16_DATA1_30), .C2(R2_n2369), .ZN(R2_n2038) );
  INV_X1 R2_U127 ( .A(R2_n2038), .ZN(R2_n417) );
  AOI222_X1 R2_U126 ( .A1(R2_n256), .A2(R2_n2386), .B1(R2_U16_DATA2_31), .B2(
        R2_n2371), .C1(R2_U16_DATA1_31), .C2(R2_n2367), .ZN(R2_n2037) );
  INV_X1 R2_U125 ( .A(R2_n2037), .ZN(R2_n418) );
  AOI222_X1 R2_U124 ( .A1(R2_n257), .A2(R2_n2389), .B1(R2_U16_DATA2_32), .B2(
        R2_n2374), .C1(R2_U16_DATA1_32), .C2(R2_n2367), .ZN(R2_n2036) );
  INV_X1 R2_U123 ( .A(R2_n2036), .ZN(R2_n419) );
  AOI222_X1 R2_U122 ( .A1(R2_n258), .A2(R2_n2386), .B1(R2_U16_DATA2_33), .B2(
        R2_n2374), .C1(R2_U16_DATA1_33), .C2(R2_n2368), .ZN(R2_n2035) );
  INV_X1 R2_U121 ( .A(R2_n2035), .ZN(R2_n420) );
  AOI222_X1 R2_U120 ( .A1(R2_n259), .A2(R2_n2390), .B1(R2_U16_DATA2_34), .B2(
        R2_n2374), .C1(R2_U16_DATA1_34), .C2(R2_n2369), .ZN(R2_n2034) );
  INV_X1 R2_U119 ( .A(R2_n2034), .ZN(R2_n421) );
  AOI222_X1 R2_U118 ( .A1(R2_n296), .A2(R2_n2387), .B1(R2_U16_DATA2_71), .B2(
        R2_n2374), .C1(R2_U16_DATA1_71), .C2(R2_n2365), .ZN(R2_n1997) );
  INV_X1 R2_U117 ( .A(R2_n1997), .ZN(R2_n458) );
  AOI222_X1 R2_U116 ( .A1(R2_n297), .A2(R2_n2387), .B1(R2_U16_DATA2_72), .B2(
        R2_n2371), .C1(R2_U16_DATA1_72), .C2(R2_n2365), .ZN(R2_n1996) );
  INV_X1 R2_U115 ( .A(R2_n1996), .ZN(R2_n459) );
  AOI222_X1 R2_U114 ( .A1(R2_n298), .A2(R2_n2387), .B1(R2_U16_DATA2_73), .B2(
        R2_n1940), .C1(R2_U16_DATA1_73), .C2(R2_n2369), .ZN(R2_n1995) );
  INV_X1 R2_U113 ( .A(R2_n1995), .ZN(R2_n460) );
  AOI222_X1 R2_U112 ( .A1(R2_n299), .A2(R2_n2387), .B1(R2_U16_DATA2_74), .B2(
        R2_n2371), .C1(R2_U16_DATA1_74), .C2(R2_n2365), .ZN(R2_n1994) );
  INV_X1 R2_U111 ( .A(R2_n1994), .ZN(R2_n461) );
  AOI222_X1 R2_U110 ( .A1(R2_n300), .A2(R2_n2387), .B1(R2_U16_DATA2_75), .B2(
        R2_n2373), .C1(R2_U16_DATA1_75), .C2(R2_n2365), .ZN(R2_n1993) );
  INV_X1 R2_U109 ( .A(R2_n1993), .ZN(R2_n462) );
  AOI222_X1 R2_U108 ( .A1(R2_n301), .A2(R2_n2387), .B1(R2_U16_DATA2_76), .B2(
        R2_n2374), .C1(R2_U16_DATA1_76), .C2(R2_n2367), .ZN(R2_n1992) );
  INV_X1 R2_U107 ( .A(R2_n1992), .ZN(R2_n463) );
  AOI222_X1 R2_U106 ( .A1(R2_n302), .A2(R2_n2387), .B1(R2_U16_DATA2_77), .B2(
        R2_n1940), .C1(R2_U16_DATA1_77), .C2(R2_n2365), .ZN(R2_n1991) );
  INV_X1 R2_U105 ( .A(R2_n1991), .ZN(R2_n464) );
  AOI222_X1 R2_U104 ( .A1(R2_n303), .A2(R2_n2387), .B1(R2_U16_DATA2_78), .B2(
        R2_n1940), .C1(R2_U16_DATA1_78), .C2(R2_n2365), .ZN(R2_n1990) );
  INV_X1 R2_U103 ( .A(R2_n1990), .ZN(R2_n465) );
  AOI222_X1 R2_U102 ( .A1(R2_n304), .A2(R2_n2387), .B1(R2_U16_DATA2_79), .B2(
        R2_n2373), .C1(R2_U16_DATA1_79), .C2(R2_n2365), .ZN(R2_n1989) );
  INV_X1 R2_U101 ( .A(R2_n1989), .ZN(R2_n466) );
  AOI222_X1 R2_U100 ( .A1(R2_n305), .A2(R2_n2387), .B1(R2_U16_DATA2_80), .B2(
        R2_n2373), .C1(R2_U16_DATA1_80), .C2(R2_n2369), .ZN(R2_n1988) );
  INV_X1 R2_U99 ( .A(R2_n1988), .ZN(R2_n467) );
  AOI222_X1 R2_U98 ( .A1(R2_n306), .A2(R2_n2387), .B1(R2_U16_DATA2_81), .B2(
        R2_n2373), .C1(R2_U16_DATA1_81), .C2(R2_n2365), .ZN(R2_n1987) );
  INV_X1 R2_U97 ( .A(R2_n1987), .ZN(R2_n468) );
  AOI222_X1 R2_U96 ( .A1(R2_n307), .A2(R2_n2387), .B1(R2_U16_DATA2_82), .B2(
        R2_n2373), .C1(R2_U16_DATA1_82), .C2(R2_n2365), .ZN(R2_n1986) );
  INV_X1 R2_U95 ( .A(R2_n1986), .ZN(R2_n469) );
  AOI222_X1 R2_U94 ( .A1(R2_n308), .A2(R2_n2388), .B1(R2_U16_DATA2_83), .B2(
        R2_n2373), .C1(R2_U16_DATA1_83), .C2(R2_n2367), .ZN(R2_n1985) );
  INV_X1 R2_U93 ( .A(R2_n1985), .ZN(R2_n470) );
  AOI222_X1 R2_U92 ( .A1(R2_n309), .A2(R2_n2388), .B1(R2_U16_DATA2_84), .B2(
        R2_n1940), .C1(R2_U16_DATA1_84), .C2(R2_n2367), .ZN(R2_n1984) );
  INV_X1 R2_U91 ( .A(R2_n1984), .ZN(R2_n471) );
  AOI222_X1 R2_U90 ( .A1(R2_n310), .A2(R2_n2388), .B1(R2_U16_DATA2_85), .B2(
        R2_n1940), .C1(R2_U16_DATA1_85), .C2(R2_n2367), .ZN(R2_n1983) );
  INV_X1 R2_U89 ( .A(R2_n1983), .ZN(R2_n472) );
  AOI222_X1 R2_U88 ( .A1(R2_n311), .A2(R2_n2388), .B1(R2_U16_DATA2_86), .B2(
        R2_n2371), .C1(R2_U16_DATA1_86), .C2(R2_n2367), .ZN(R2_n1982) );
  INV_X1 R2_U87 ( .A(R2_n1982), .ZN(R2_n473) );
  AOI222_X1 R2_U86 ( .A1(R2_n312), .A2(R2_n2388), .B1(R2_U16_DATA2_87), .B2(
        R2_n2370), .C1(R2_U16_DATA1_87), .C2(R2_n2367), .ZN(R2_n1981) );
  INV_X1 R2_U85 ( .A(R2_n1981), .ZN(R2_n474) );
  AOI222_X1 R2_U84 ( .A1(R2_n313), .A2(R2_n2388), .B1(R2_U16_DATA2_88), .B2(
        R2_n2371), .C1(R2_U16_DATA1_88), .C2(R2_n2367), .ZN(R2_n1980) );
  INV_X1 R2_U83 ( .A(R2_n1980), .ZN(R2_n475) );
  AOI222_X1 R2_U82 ( .A1(R2_n314), .A2(R2_n2388), .B1(R2_U16_DATA2_89), .B2(
        R2_n2373), .C1(R2_U16_DATA1_89), .C2(R2_n2367), .ZN(R2_n1979) );
  INV_X1 R2_U81 ( .A(R2_n1979), .ZN(R2_n476) );
  AOI222_X1 R2_U80 ( .A1(R2_n315), .A2(R2_n2388), .B1(R2_U16_DATA2_90), .B2(
        R2_n2371), .C1(R2_U16_DATA1_90), .C2(R2_n2367), .ZN(R2_n1978) );
  INV_X1 R2_U79 ( .A(R2_n1978), .ZN(R2_n477) );
  AOI222_X1 R2_U78 ( .A1(R2_n316), .A2(R2_n2388), .B1(R2_U16_DATA2_91), .B2(
        R2_n2373), .C1(R2_U16_DATA1_91), .C2(R2_n2367), .ZN(R2_n1977) );
  INV_X1 R2_U77 ( .A(R2_n1977), .ZN(R2_n478) );
  AOI222_X1 R2_U76 ( .A1(R2_n317), .A2(R2_n2388), .B1(R2_U16_DATA2_92), .B2(
        R2_n2373), .C1(R2_U16_DATA1_92), .C2(R2_n2367), .ZN(R2_n1976) );
  INV_X1 R2_U75 ( .A(R2_n1976), .ZN(R2_n479) );
  AOI222_X1 R2_U74 ( .A1(R2_n318), .A2(R2_n2388), .B1(R2_U16_DATA2_93), .B2(
        R2_n1940), .C1(R2_U16_DATA1_93), .C2(R2_n2367), .ZN(R2_n1975) );
  INV_X1 R2_U73 ( .A(R2_n1975), .ZN(R2_n480) );
  AOI222_X1 R2_U72 ( .A1(R2_n319), .A2(R2_n2388), .B1(R2_U16_DATA2_94), .B2(
        R2_n2370), .C1(R2_U16_DATA1_94), .C2(R2_n2367), .ZN(R2_n1974) );
  INV_X1 R2_U71 ( .A(R2_n1974), .ZN(R2_n481) );
  NOR2_X1 R2_U70 ( .A1(n3261), .A2(R2_n2348), .ZN(R2_n2332) );
  NAND2_X1 R2_U69 ( .A1(R2_n2337), .A2(R2_r332_A_1_), .ZN(R2_n2335) );
  OAI21_X1 R2_U68 ( .B1(R2_n1806), .B2(R2_n2328), .A(R2_n2329), .ZN(R2_n2338)
         );
  OAI22_X1 R2_U67 ( .A1(R2_n1), .A2(R2_n1805), .B1(R2_r332_A_1_), .B2(R2_n2330), .ZN(R2_n2339) );
  OAI22_X1 R2_U66 ( .A1(R2_n1), .A2(R2_n1804), .B1(R2_n1805), .B2(R2_n2330), 
        .ZN(R2_n2340) );
  OAI21_X1 R2_U65 ( .B1(n3261), .B2(R2_r332_A_0_), .A(R2_n2328), .ZN(R2_n2331)
         );
  NOR2_X1 R2_U63 ( .A1(n3261), .A2(R2_n1514), .ZN(R2_n2334) );
  NOR3_X1 R2_U62 ( .A1(R2_r332_A_2_), .A2(R2_r332_A_3_), .A3(R2_r332_A_0_), 
        .ZN(R2_n2337) );
  INV_X1 R2_U59 ( .A(R2_n2331), .ZN(R2_n1) );
  INV_X1 R2_U58 ( .A(R2_n2334), .ZN(R2_n1808) );
  NOR2_X1 R2_U57 ( .A1(R2_n1808), .A2(R2_n2335), .ZN(R2_n2069) );
  BUF_X1 R2_U56 ( .A(R2_n2366), .Z(R2_n2368) );
  INV_X1 R2_U55 ( .A(R2_n2069), .ZN(R2_n1802) );
  BUF_X1 R2_U51 ( .A(R2_n2354), .Z(R2_n2364) );
  BUF_X1 R2_U50 ( .A(R2_n2354), .Z(R2_n2362) );
  INV_X1 R2_U48 ( .A(R2_n2343), .ZN(R2_n2344) );
  INV_X1 R2_U47 ( .A(R2_n2343), .ZN(R2_n2345) );
  INV_X1 R2_U46 ( .A(R2_n2343), .ZN(R2_n2346) );
  INV_X1 R2_U45 ( .A(R2_n2343), .ZN(R2_n2349) );
  INV_X1 R2_U44 ( .A(R2_n2343), .ZN(R2_n2347) );
  INV_X1 R2_U43 ( .A(R2_n2200), .ZN(R2_n2348) );
  INV_X1 R2_U41 ( .A(R2_n1811), .ZN(R2_n2382) );
  INV_X1 R2_U40 ( .A(R2_n1811), .ZN(R2_n2381) );
  INV_X1 R2_U39 ( .A(R2_n1811), .ZN(R2_n2378) );
  INV_X1 R2_U38 ( .A(R2_n2376), .ZN(R2_n2377) );
  INV_X1 R2_U37 ( .A(R2_n2376), .ZN(R2_n2380) );
  INV_X1 R2_U36 ( .A(R2_n1811), .ZN(R2_n2379) );
  INV_X1 R2_U35 ( .A(R2_n2071), .ZN(R2_n2356) );
  INV_X1 R2_U34 ( .A(R2_n2071), .ZN(R2_n2355) );
  INV_X1 R2_U33 ( .A(R2_n2071), .ZN(R2_n2360) );
  INV_X1 R2_U32 ( .A(R2_n2071), .ZN(R2_n2359) );
  INV_X1 R2_U31 ( .A(R2_n2071), .ZN(R2_n2358) );
  INV_X1 R2_U30 ( .A(R2_n2071), .ZN(R2_n2357) );
  CLKBUF_X1 R2_U29 ( .A(R2_n2354), .Z(R2_n2363) );
  CLKBUF_X1 R2_U28 ( .A(R2_n2071), .Z(R2_n2354) );
  CLKBUF_X1 R2_U27 ( .A(R2_n2375), .Z(R2_n2385) );
  CLKBUF_X1 R2_U26 ( .A(R2_n2375), .Z(R2_n2384) );
  CLKBUF_X1 R2_U25 ( .A(R2_n2375), .Z(R2_n2383) );
  CLKBUF_X1 R2_U22 ( .A(R2_n2352), .Z(R2_n2351) );
  CLKBUF_X1 R2_U21 ( .A(R2_n2200), .Z(R2_n2350) );
  CLKBUF_X1 R2_U19 ( .A(R2_n2343), .Z(R2_n2352) );
  CLKBUF_X1 R2_U16 ( .A(R2_n1940), .Z(R2_n2370) );
  CLKBUF_X1 R2_U15 ( .A(R2_n1940), .Z(R2_n2371) );
  CLKBUF_X1 R2_U13 ( .A(R2_n2370), .Z(R2_n2372) );
  CLKBUF_X1 R2_U11 ( .A(R2_n2366), .Z(R2_n2367) );
  CLKBUF_X1 R2_U10 ( .A(R2_n2366), .Z(R2_n2369) );
  CLKBUF_X1 R2_U9 ( .A(R2_n1941), .Z(R2_n2366) );
  NAND4_X1 R2_U1060 ( .A1(R2_n2376), .A2(R2_n2390), .A3(R2_n2332), .A4(
        R2_n2071), .ZN(R2_n2328) );
  NAND3_X1 R2_U1059 ( .A1(R2_n2328), .A2(R2_n1809), .A3(R2_r332_A_0_), .ZN(
        R2_n2330) );
  NAND3_X1 R2_U1058 ( .A1(R2_n1806), .A2(R2_n1809), .A3(R2_n2328), .ZN(
        R2_n2329) );
  DFF_X1 R2_temp_add_data_reg_127_ ( .D(R2_n1800), .CK(clk), .Q(n3390) );
  DFF_X1 R2_temp_add_data_reg_126_ ( .D(R2_n1799), .CK(clk), .Q(n3389) );
  DFF_X1 R2_temp_add_data_reg_125_ ( .D(R2_n1798), .CK(clk), .Q(n3388) );
  DFF_X1 R2_temp_add_data_reg_124_ ( .D(R2_n1797), .CK(clk), .Q(n3387) );
  DFF_X1 R2_temp_add_data_reg_123_ ( .D(R2_n1796), .CK(clk), .Q(n3386) );
  DFF_X1 R2_temp_add_data_reg_122_ ( .D(R2_n1795), .CK(clk), .Q(n3385) );
  DFF_X1 R2_temp_add_data_reg_121_ ( .D(R2_n1794), .CK(clk), .Q(n3384) );
  DFF_X1 R2_temp_add_data_reg_120_ ( .D(R2_n1793), .CK(clk), .Q(n3383) );
  DFF_X1 R2_temp_add_data_reg_119_ ( .D(R2_n1792), .CK(clk), .Q(n3382) );
  DFF_X1 R2_temp_add_data_reg_118_ ( .D(R2_n1791), .CK(clk), .Q(n3381) );
  DFF_X1 R2_temp_add_data_reg_117_ ( .D(R2_n1790), .CK(clk), .Q(n3380) );
  DFF_X1 R2_temp_add_data_reg_116_ ( .D(R2_n1789), .CK(clk), .Q(n3379) );
  DFF_X1 R2_temp_add_data_reg_115_ ( .D(R2_n1788), .CK(clk), .Q(n3378) );
  DFF_X1 R2_temp_add_data_reg_114_ ( .D(R2_n1787), .CK(clk), .Q(n3377) );
  DFF_X1 R2_temp_add_data_reg_113_ ( .D(R2_n1786), .CK(clk), .Q(n3376) );
  DFF_X1 R2_temp_add_data_reg_112_ ( .D(R2_n1785), .CK(clk), .Q(n3375) );
  DFF_X1 R2_temp_add_data_reg_111_ ( .D(R2_n1784), .CK(clk), .Q(n3374) );
  DFF_X1 R2_temp_add_data_reg_110_ ( .D(R2_n1783), .CK(clk), .Q(n3373) );
  DFF_X1 R2_temp_add_data_reg_109_ ( .D(R2_n1782), .CK(clk), .Q(n3372) );
  DFF_X1 R2_temp_add_data_reg_108_ ( .D(R2_n1781), .CK(clk), .Q(n3371) );
  DFF_X1 R2_temp_add_data_reg_107_ ( .D(R2_n1780), .CK(clk), .Q(n3370) );
  DFF_X1 R2_temp_add_data_reg_106_ ( .D(R2_n1779), .CK(clk), .Q(n3369) );
  DFF_X1 R2_temp_add_data_reg_105_ ( .D(R2_n1778), .CK(clk), .Q(n3368) );
  DFF_X1 R2_temp_add_data_reg_104_ ( .D(R2_n1777), .CK(clk), .Q(n3367) );
  DFF_X1 R2_temp_add_data_reg_103_ ( .D(R2_n1776), .CK(clk), .Q(n3366) );
  DFF_X1 R2_temp_add_data_reg_102_ ( .D(R2_n1775), .CK(clk), .Q(n3365) );
  DFF_X1 R2_temp_add_data_reg_101_ ( .D(R2_n1774), .CK(clk), .Q(n3364) );
  DFF_X1 R2_temp_add_data_reg_100_ ( .D(R2_n1773), .CK(clk), .Q(n3363) );
  DFF_X1 R2_temp_add_data_reg_99_ ( .D(R2_n1772), .CK(clk), .Q(n3362) );
  DFF_X1 R2_temp_add_data_reg_98_ ( .D(R2_n1128), .CK(clk), .Q(n3361) );
  DFF_X1 R2_temp_add_data_reg_97_ ( .D(R2_n1127), .CK(clk), .Q(n3360) );
  DFF_X1 R2_temp_add_data_reg_96_ ( .D(R2_n1126), .CK(clk), .Q(n3359) );
  DFF_X1 R2_temp_add_data_reg_95_ ( .D(R2_n1125), .CK(clk), .Q(n3358) );
  DFF_X1 R2_temp_add_data_reg_94_ ( .D(R2_n1124), .CK(clk), .Q(n3357) );
  DFF_X1 R2_temp_add_data_reg_93_ ( .D(R2_n1123), .CK(clk), .Q(n3356) );
  DFF_X1 R2_temp_add_data_reg_92_ ( .D(R2_n1122), .CK(clk), .Q(n3355) );
  DFF_X1 R2_temp_add_data_reg_91_ ( .D(R2_n1121), .CK(clk), .Q(n3354) );
  DFF_X1 R2_temp_add_data_reg_90_ ( .D(R2_n1120), .CK(clk), .Q(n3353) );
  DFF_X1 R2_temp_add_data_reg_89_ ( .D(R2_n1119), .CK(clk), .Q(n3352) );
  DFF_X1 R2_temp_add_data_reg_88_ ( .D(R2_n1118), .CK(clk), .Q(n3351) );
  DFF_X1 R2_temp_add_data_reg_87_ ( .D(R2_n1117), .CK(clk), .Q(n3350) );
  DFF_X1 R2_temp_add_data_reg_86_ ( .D(R2_n1116), .CK(clk), .Q(n3349) );
  DFF_X1 R2_temp_add_data_reg_85_ ( .D(R2_n1115), .CK(clk), .Q(n3348) );
  DFF_X1 R2_temp_add_data_reg_84_ ( .D(R2_n1114), .CK(clk), .Q(n3347) );
  DFF_X1 R2_temp_add_data_reg_83_ ( .D(R2_n1113), .CK(clk), .Q(n3346) );
  DFF_X1 R2_temp_add_data_reg_82_ ( .D(R2_n1112), .CK(clk), .Q(n3345) );
  DFF_X1 R2_temp_add_data_reg_81_ ( .D(R2_n1111), .CK(clk), .Q(n3344) );
  DFF_X1 R2_temp_add_data_reg_80_ ( .D(R2_n1110), .CK(clk), .Q(n3343) );
  DFF_X1 R2_temp_add_data_reg_79_ ( .D(R2_n1109), .CK(clk), .Q(n3342) );
  DFF_X1 R2_temp_add_data_reg_78_ ( .D(R2_n1108), .CK(clk), .Q(n3341) );
  DFF_X1 R2_temp_add_data_reg_77_ ( .D(R2_n1107), .CK(clk), .Q(n3340) );
  DFF_X1 R2_temp_add_data_reg_76_ ( .D(R2_n1106), .CK(clk), .Q(n3339) );
  DFF_X1 R2_temp_add_data_reg_75_ ( .D(R2_n1105), .CK(clk), .Q(n3338) );
  DFF_X1 R2_temp_add_data_reg_74_ ( .D(R2_n1104), .CK(clk), .Q(n3337) );
  DFF_X1 R2_temp_add_data_reg_73_ ( .D(R2_n1103), .CK(clk), .Q(n3336) );
  DFF_X1 R2_temp_add_data_reg_72_ ( .D(R2_n1102), .CK(clk), .Q(n3335) );
  DFF_X1 R2_temp_add_data_reg_71_ ( .D(R2_n1101), .CK(clk), .Q(n3334) );
  DFF_X1 R2_temp_add_data_reg_70_ ( .D(R2_n1100), .CK(clk), .Q(n3333) );
  DFF_X1 R2_temp_add_data_reg_69_ ( .D(R2_n1099), .CK(clk), .Q(n3332) );
  DFF_X1 R2_temp_add_data_reg_68_ ( .D(R2_n1098), .CK(clk), .Q(n3331) );
  DFF_X1 R2_temp_add_data_reg_67_ ( .D(R2_n1097), .CK(clk), .Q(n3330) );
  DFF_X1 R2_temp_add_data_reg_66_ ( .D(R2_n1096), .CK(clk), .Q(n3329) );
  DFF_X1 R2_temp_add_data_reg_65_ ( .D(R2_n1095), .CK(clk), .Q(n3328) );
  DFF_X1 R2_temp_add_data_reg_64_ ( .D(R2_n1094), .CK(clk), .Q(n3327) );
  DFF_X1 R2_temp_add_data_reg_63_ ( .D(R2_n1093), .CK(clk), .Q(n3326) );
  DFF_X1 R2_temp_add_data_reg_62_ ( .D(R2_n1092), .CK(clk), .Q(n3325) );
  DFF_X1 R2_temp_add_data_reg_61_ ( .D(R2_n1091), .CK(clk), .Q(n3324) );
  DFF_X1 R2_temp_add_data_reg_60_ ( .D(R2_n1090), .CK(clk), .Q(n3323) );
  DFF_X1 R2_temp_add_data_reg_59_ ( .D(R2_n1089), .CK(clk), .Q(n3322) );
  DFF_X1 R2_temp_add_data_reg_58_ ( .D(R2_n1088), .CK(clk), .Q(n3321) );
  DFF_X1 R2_temp_add_data_reg_57_ ( .D(R2_n1087), .CK(clk), .Q(n3320) );
  DFF_X1 R2_temp_add_data_reg_56_ ( .D(R2_n1086), .CK(clk), .Q(n3319) );
  DFF_X1 R2_temp_add_data_reg_55_ ( .D(R2_n1085), .CK(clk), .Q(n3318) );
  DFF_X1 R2_temp_add_data_reg_54_ ( .D(R2_n1084), .CK(clk), .Q(n3317) );
  DFF_X1 R2_temp_add_data_reg_53_ ( .D(R2_n1083), .CK(clk), .Q(n3316) );
  DFF_X1 R2_temp_add_data_reg_52_ ( .D(R2_n1082), .CK(clk), .Q(n3315) );
  DFF_X1 R2_temp_add_data_reg_51_ ( .D(R2_n1081), .CK(clk), .Q(n3314) );
  DFF_X1 R2_temp_add_data_reg_50_ ( .D(R2_n1080), .CK(clk), .Q(n3313) );
  DFF_X1 R2_temp_add_data_reg_49_ ( .D(R2_n1079), .CK(clk), .Q(n3312) );
  DFF_X1 R2_temp_add_data_reg_48_ ( .D(R2_n1078), .CK(clk), .Q(n3311) );
  DFF_X1 R2_temp_add_data_reg_47_ ( .D(R2_n1077), .CK(clk), .Q(n3310) );
  DFF_X1 R2_temp_add_data_reg_46_ ( .D(R2_n1076), .CK(clk), .Q(n3309) );
  DFF_X1 R2_temp_add_data_reg_45_ ( .D(R2_n1075), .CK(clk), .Q(n3308) );
  DFF_X1 R2_temp_add_data_reg_44_ ( .D(R2_n1074), .CK(clk), .Q(n3307) );
  DFF_X1 R2_temp_add_data_reg_43_ ( .D(R2_n1073), .CK(clk), .Q(n3306) );
  DFF_X1 R2_temp_add_data_reg_42_ ( .D(R2_n1072), .CK(clk), .Q(n3305) );
  DFF_X1 R2_temp_add_data_reg_41_ ( .D(R2_n1071), .CK(clk), .Q(n3304) );
  DFF_X1 R2_temp_add_data_reg_40_ ( .D(R2_n1070), .CK(clk), .Q(n3303) );
  DFF_X1 R2_temp_add_data_reg_39_ ( .D(R2_n1069), .CK(clk), .Q(n3302) );
  DFF_X1 R2_temp_add_data_reg_38_ ( .D(R2_n1068), .CK(clk), .Q(n3301) );
  DFF_X1 R2_temp_add_data_reg_37_ ( .D(R2_n1067), .CK(clk), .Q(n3300) );
  DFF_X1 R2_temp_add_data_reg_36_ ( .D(R2_n1066), .CK(clk), .Q(n3299) );
  DFF_X1 R2_temp_add_data_reg_35_ ( .D(R2_n1065), .CK(clk), .Q(n3298) );
  DFF_X1 R2_temp_add_data_reg_34_ ( .D(R2_n1064), .CK(clk), .Q(n3297) );
  DFF_X1 R2_temp_add_data_reg_33_ ( .D(R2_n1063), .CK(clk), .Q(n3296) );
  DFF_X1 R2_temp_add_data_reg_32_ ( .D(R2_n1062), .CK(clk), .Q(n3295) );
  DFF_X1 R2_temp_add_data_reg_31_ ( .D(R2_n1061), .CK(clk), .Q(n3294) );
  DFF_X1 R2_temp_add_data_reg_30_ ( .D(R2_n1060), .CK(clk), .Q(n3293) );
  DFF_X1 R2_temp_add_data_reg_29_ ( .D(R2_n1059), .CK(clk), .Q(n3292) );
  DFF_X1 R2_temp_add_data_reg_28_ ( .D(R2_n1058), .CK(clk), .Q(n3291) );
  DFF_X1 R2_temp_add_data_reg_27_ ( .D(R2_n1057), .CK(clk), .Q(n3290) );
  DFF_X1 R2_temp_add_data_reg_26_ ( .D(R2_n1056), .CK(clk), .Q(n3289) );
  DFF_X1 R2_temp_add_data_reg_25_ ( .D(R2_n1055), .CK(clk), .Q(n3288) );
  DFF_X1 R2_temp_add_data_reg_24_ ( .D(R2_n1054), .CK(clk), .Q(n3287) );
  DFF_X1 R2_temp_add_data_reg_23_ ( .D(R2_n1053), .CK(clk), .Q(n3286) );
  DFF_X1 R2_temp_add_data_reg_22_ ( .D(R2_n1052), .CK(clk), .Q(n3285) );
  DFF_X1 R2_temp_add_data_reg_21_ ( .D(R2_n1051), .CK(clk), .Q(n3284) );
  DFF_X1 R2_temp_add_data_reg_20_ ( .D(R2_n1050), .CK(clk), .Q(n3283) );
  DFF_X1 R2_temp_add_data_reg_19_ ( .D(R2_n1049), .CK(clk), .Q(n3282) );
  DFF_X1 R2_temp_add_data_reg_18_ ( .D(R2_n1048), .CK(clk), .Q(n3281) );
  DFF_X1 R2_temp_add_data_reg_17_ ( .D(R2_n1047), .CK(clk), .Q(n3280) );
  DFF_X1 R2_temp_add_data_reg_16_ ( .D(R2_n1046), .CK(clk), .Q(n3279) );
  DFF_X1 R2_temp_add_data_reg_15_ ( .D(R2_n1045), .CK(clk), .Q(n3278) );
  DFF_X1 R2_temp_add_data_reg_14_ ( .D(R2_n1044), .CK(clk), .Q(n3277) );
  DFF_X1 R2_temp_add_data_reg_13_ ( .D(R2_n1043), .CK(clk), .Q(n3276) );
  DFF_X1 R2_temp_add_data_reg_12_ ( .D(R2_n1042), .CK(clk), .Q(n3275) );
  DFF_X1 R2_temp_add_data_reg_11_ ( .D(R2_n1041), .CK(clk), .Q(n3274) );
  DFF_X1 R2_temp_add_data_reg_10_ ( .D(R2_n1040), .CK(clk), .Q(n3273) );
  DFF_X1 R2_temp_add_data_reg_9_ ( .D(R2_n1039), .CK(clk), .Q(n3272) );
  DFF_X1 R2_temp_add_data_reg_8_ ( .D(R2_n1038), .CK(clk), .Q(n3271) );
  DFF_X1 R2_temp_add_data_reg_7_ ( .D(R2_n1037), .CK(clk), .Q(n3270) );
  DFF_X1 R2_temp_add_data_reg_6_ ( .D(R2_n1036), .CK(clk), .Q(n3269) );
  DFF_X1 R2_temp_add_data_reg_5_ ( .D(R2_n1035), .CK(clk), .Q(n3268) );
  DFF_X1 R2_temp_add_data_reg_4_ ( .D(R2_n1034), .CK(clk), .Q(n3267) );
  DFF_X1 R2_temp_add_data_reg_3_ ( .D(R2_n1033), .CK(clk), .Q(n3266) );
  DFF_X1 R2_temp_add_data_reg_2_ ( .D(R2_n1032), .CK(clk), .Q(n3265) );
  DFF_X1 R2_temp_add_data_reg_1_ ( .D(R2_n1031), .CK(clk), .Q(n3264) );
  DFF_X1 R2_temp_add_data_reg_0_ ( .D(R2_n1030), .CK(clk), .Q(n3263) );
  DLH_X1 R2_add_in_data_reg_127_ ( .G(R2_n2402), .D(R2_n352), .Q(R2_n999) );
  DFF_X1 R2_temp_mix_data_reg_127_ ( .D(R2_n1029), .CK(clk), .Q(R2_n352) );
  DLH_X1 R2_add_in_data_reg_126_ ( .G(R2_n2403), .D(R2_n351), .Q(R2_n998) );
  DFF_X1 R2_temp_mix_data_reg_126_ ( .D(R2_n1028), .CK(clk), .Q(R2_n351) );
  DLH_X1 R2_add_in_data_reg_125_ ( .G(R2_n2404), .D(R2_n350), .Q(R2_n997) );
  DFF_X1 R2_temp_mix_data_reg_125_ ( .D(R2_n1027), .CK(clk), .Q(R2_n350) );
  DLH_X1 R2_add_in_data_reg_124_ ( .G(R2_U23_Z_1), .D(R2_n349), .Q(R2_n996) );
  DFF_X1 R2_temp_mix_data_reg_124_ ( .D(R2_n1026), .CK(clk), .Q(R2_n349) );
  DLH_X1 R2_add_in_data_reg_123_ ( .G(R2_n2401), .D(R2_n348), .Q(R2_n995) );
  DFF_X1 R2_temp_mix_data_reg_123_ ( .D(R2_n1025), .CK(clk), .Q(R2_n348) );
  DLH_X1 R2_add_in_data_reg_122_ ( .G(R2_U23_Z_1), .D(R2_n347), .Q(R2_n994) );
  DFF_X1 R2_temp_mix_data_reg_122_ ( .D(R2_n1024), .CK(clk), .Q(R2_n347) );
  DLH_X1 R2_add_in_data_reg_121_ ( .G(R2_n2403), .D(R2_n346), .Q(R2_n993) );
  DFF_X1 R2_temp_mix_data_reg_121_ ( .D(R2_n1023), .CK(clk), .Q(R2_n346) );
  DLH_X1 R2_add_in_data_reg_120_ ( .G(R2_n2398), .D(R2_n345), .Q(R2_n992) );
  DFF_X1 R2_temp_mix_data_reg_120_ ( .D(R2_n1022), .CK(clk), .Q(R2_n345) );
  DLH_X1 R2_add_in_data_reg_119_ ( .G(R2_U23_Z_1), .D(R2_n344), .Q(R2_n991) );
  DFF_X1 R2_temp_mix_data_reg_119_ ( .D(R2_n1021), .CK(clk), .Q(R2_n344) );
  DLH_X1 R2_add_in_data_reg_118_ ( .G(R2_n2398), .D(R2_n343), .Q(R2_n990) );
  DFF_X1 R2_temp_mix_data_reg_118_ ( .D(R2_n1020), .CK(clk), .Q(R2_n343) );
  DLH_X1 R2_add_in_data_reg_117_ ( .G(R2_U23_Z_1), .D(R2_n342), .Q(R2_n989) );
  DFF_X1 R2_temp_mix_data_reg_117_ ( .D(R2_n1019), .CK(clk), .Q(R2_n342) );
  DLH_X1 R2_add_in_data_reg_116_ ( .G(R2_n2404), .D(R2_n341), .Q(R2_n988) );
  DFF_X1 R2_temp_mix_data_reg_116_ ( .D(R2_n1018), .CK(clk), .Q(R2_n341) );
  DLH_X1 R2_add_in_data_reg_115_ ( .G(R2_n2400), .D(R2_n340), .Q(R2_n987) );
  DFF_X1 R2_temp_mix_data_reg_115_ ( .D(R2_n1017), .CK(clk), .Q(R2_n340) );
  DLH_X1 R2_add_in_data_reg_114_ ( .G(R2_n2404), .D(R2_n339), .Q(R2_n986) );
  DFF_X1 R2_temp_mix_data_reg_114_ ( .D(R2_n1016), .CK(clk), .Q(R2_n339) );
  DLH_X1 R2_add_in_data_reg_113_ ( .G(R2_n2404), .D(R2_n338), .Q(R2_n985) );
  DFF_X1 R2_temp_mix_data_reg_113_ ( .D(R2_n1015), .CK(clk), .Q(R2_n338) );
  DLH_X1 R2_add_in_data_reg_112_ ( .G(R2_n2399), .D(R2_n337), .Q(R2_n984) );
  DFF_X1 R2_temp_mix_data_reg_112_ ( .D(R2_n1014), .CK(clk), .Q(R2_n337) );
  DLH_X1 R2_add_in_data_reg_111_ ( .G(R2_n2400), .D(R2_n336), .Q(R2_n983) );
  DFF_X1 R2_temp_mix_data_reg_111_ ( .D(R2_n1013), .CK(clk), .Q(R2_n336) );
  DLH_X1 R2_add_in_data_reg_110_ ( .G(R2_n2398), .D(R2_n335), .Q(R2_n982) );
  DFF_X1 R2_temp_mix_data_reg_110_ ( .D(R2_n1012), .CK(clk), .Q(R2_n335) );
  DLH_X1 R2_add_in_data_reg_109_ ( .G(R2_n2402), .D(R2_n334), .Q(R2_n981) );
  DFF_X1 R2_temp_mix_data_reg_109_ ( .D(R2_n1011), .CK(clk), .Q(R2_n334) );
  DLH_X1 R2_add_in_data_reg_108_ ( .G(R2_n2399), .D(R2_n333), .Q(R2_n980) );
  DFF_X1 R2_temp_mix_data_reg_108_ ( .D(R2_n1010), .CK(clk), .Q(R2_n333) );
  DLH_X1 R2_add_in_data_reg_107_ ( .G(R2_n2398), .D(R2_n332), .Q(R2_n979) );
  DFF_X1 R2_temp_mix_data_reg_107_ ( .D(R2_n1009), .CK(clk), .Q(R2_n332) );
  DLH_X1 R2_add_in_data_reg_106_ ( .G(R2_n2399), .D(R2_n331), .Q(R2_n978) );
  DFF_X1 R2_temp_mix_data_reg_106_ ( .D(R2_n1008), .CK(clk), .Q(R2_n331) );
  DLH_X1 R2_add_in_data_reg_105_ ( .G(R2_n2404), .D(R2_n330), .Q(R2_n977) );
  DFF_X1 R2_temp_mix_data_reg_105_ ( .D(R2_n1007), .CK(clk), .Q(R2_n330) );
  DLH_X1 R2_add_in_data_reg_104_ ( .G(R2_n2402), .D(R2_n329), .Q(R2_n976) );
  DFF_X1 R2_temp_mix_data_reg_104_ ( .D(R2_n1006), .CK(clk), .Q(R2_n329) );
  DLH_X1 R2_add_in_data_reg_103_ ( .G(R2_n2398), .D(R2_n328), .Q(R2_n975) );
  DFF_X1 R2_temp_mix_data_reg_103_ ( .D(R2_n1005), .CK(clk), .Q(R2_n328) );
  DLH_X1 R2_add_in_data_reg_102_ ( .G(R2_U23_Z_1), .D(R2_n327), .Q(R2_n974) );
  DFF_X1 R2_temp_mix_data_reg_102_ ( .D(R2_n1004), .CK(clk), .Q(R2_n327) );
  DLH_X1 R2_add_in_data_reg_101_ ( .G(R2_n2402), .D(R2_n326), .Q(R2_n973) );
  DFF_X1 R2_temp_mix_data_reg_101_ ( .D(R2_n1003), .CK(clk), .Q(R2_n326) );
  DLH_X1 R2_add_in_data_reg_100_ ( .G(R2_n2401), .D(R2_n325), .Q(R2_n972) );
  DFF_X1 R2_temp_mix_data_reg_100_ ( .D(R2_n1002), .CK(clk), .Q(R2_n325) );
  DLH_X1 R2_add_in_data_reg_99_ ( .G(R2_U23_Z_1), .D(R2_n324), .Q(R2_n971) );
  DFF_X1 R2_temp_mix_data_reg_99_ ( .D(R2_n1001), .CK(clk), .Q(R2_n324) );
  DLH_X1 R2_add_in_data_reg_98_ ( .G(R2_n2404), .D(R2_n323), .Q(R2_n970) );
  DFF_X1 R2_temp_mix_data_reg_98_ ( .D(R2_n614), .CK(clk), .Q(R2_n323) );
  DLH_X1 R2_add_in_data_reg_97_ ( .G(R2_U23_Z_1), .D(R2_n322), .Q(R2_n969) );
  DFF_X1 R2_temp_mix_data_reg_97_ ( .D(R2_n613), .CK(clk), .Q(R2_n322) );
  DLH_X1 R2_add_in_data_reg_96_ ( .G(R2_U23_Z_1), .D(R2_n321), .Q(R2_n968) );
  DFF_X1 R2_temp_mix_data_reg_96_ ( .D(R2_n612), .CK(clk), .Q(R2_n321) );
  DLH_X1 R2_add_in_data_reg_95_ ( .G(R2_n2401), .D(R2_n320), .Q(R2_n967) );
  DFF_X1 R2_temp_mix_data_reg_95_ ( .D(R2_n611), .CK(clk), .Q(R2_n320) );
  DLH_X1 R2_add_in_data_reg_94_ ( .G(R2_n2399), .D(R2_n319), .Q(R2_n966) );
  DFF_X1 R2_temp_mix_data_reg_94_ ( .D(R2_n481), .CK(clk), .Q(R2_n319) );
  DLH_X1 R2_add_in_data_reg_93_ ( .G(R2_n2400), .D(R2_n318), .Q(R2_n965) );
  DFF_X1 R2_temp_mix_data_reg_93_ ( .D(R2_n480), .CK(clk), .Q(R2_n318) );
  DLH_X1 R2_add_in_data_reg_92_ ( .G(R2_n2403), .D(R2_n317), .Q(R2_n964) );
  DFF_X1 R2_temp_mix_data_reg_92_ ( .D(R2_n479), .CK(clk), .Q(R2_n317) );
  DLH_X1 R2_add_in_data_reg_91_ ( .G(R2_n2399), .D(R2_n316), .Q(R2_n963) );
  DFF_X1 R2_temp_mix_data_reg_91_ ( .D(R2_n478), .CK(clk), .Q(R2_n316) );
  DLH_X1 R2_add_in_data_reg_90_ ( .G(R2_n2404), .D(R2_n315), .Q(R2_n962) );
  DFF_X1 R2_temp_mix_data_reg_90_ ( .D(R2_n477), .CK(clk), .Q(R2_n315) );
  DLH_X1 R2_add_in_data_reg_89_ ( .G(R2_U23_Z_1), .D(R2_n314), .Q(R2_n961) );
  DFF_X1 R2_temp_mix_data_reg_89_ ( .D(R2_n476), .CK(clk), .Q(R2_n314) );
  DLH_X1 R2_add_in_data_reg_88_ ( .G(R2_n2398), .D(R2_n313), .Q(R2_n960) );
  DFF_X1 R2_temp_mix_data_reg_88_ ( .D(R2_n475), .CK(clk), .Q(R2_n313) );
  DLH_X1 R2_add_in_data_reg_87_ ( .G(R2_n2398), .D(R2_n312), .Q(R2_n959) );
  DFF_X1 R2_temp_mix_data_reg_87_ ( .D(R2_n474), .CK(clk), .Q(R2_n312) );
  DLH_X1 R2_add_in_data_reg_86_ ( .G(R2_n2398), .D(R2_n311), .Q(R2_n958) );
  DFF_X1 R2_temp_mix_data_reg_86_ ( .D(R2_n473), .CK(clk), .Q(R2_n311) );
  DLH_X1 R2_add_in_data_reg_85_ ( .G(R2_n2398), .D(R2_n310), .Q(R2_n957) );
  DFF_X1 R2_temp_mix_data_reg_85_ ( .D(R2_n472), .CK(clk), .Q(R2_n310) );
  DLH_X1 R2_add_in_data_reg_84_ ( .G(R2_U23_Z_1), .D(R2_n309), .Q(R2_n956) );
  DFF_X1 R2_temp_mix_data_reg_84_ ( .D(R2_n471), .CK(clk), .Q(R2_n309) );
  DLH_X1 R2_add_in_data_reg_83_ ( .G(R2_n2398), .D(R2_n308), .Q(R2_n955) );
  DFF_X1 R2_temp_mix_data_reg_83_ ( .D(R2_n470), .CK(clk), .Q(R2_n308) );
  DLH_X1 R2_add_in_data_reg_82_ ( .G(R2_n2398), .D(R2_n307), .Q(R2_n954) );
  DFF_X1 R2_temp_mix_data_reg_82_ ( .D(R2_n469), .CK(clk), .Q(R2_n307) );
  DLH_X1 R2_add_in_data_reg_81_ ( .G(R2_n2401), .D(R2_n306), .Q(R2_n953) );
  DFF_X1 R2_temp_mix_data_reg_81_ ( .D(R2_n468), .CK(clk), .Q(R2_n306) );
  DLH_X1 R2_add_in_data_reg_80_ ( .G(R2_n2399), .D(R2_n305), .Q(R2_n952) );
  DFF_X1 R2_temp_mix_data_reg_80_ ( .D(R2_n467), .CK(clk), .Q(R2_n305) );
  DLH_X1 R2_add_in_data_reg_79_ ( .G(R2_n2403), .D(R2_n304), .Q(R2_n951) );
  DFF_X1 R2_temp_mix_data_reg_79_ ( .D(R2_n466), .CK(clk), .Q(R2_n304) );
  DLH_X1 R2_add_in_data_reg_78_ ( .G(R2_U23_Z_1), .D(R2_n303), .Q(R2_n950) );
  DFF_X1 R2_temp_mix_data_reg_78_ ( .D(R2_n465), .CK(clk), .Q(R2_n303) );
  DLH_X1 R2_add_in_data_reg_77_ ( .G(R2_n2401), .D(R2_n302), .Q(R2_n949) );
  DFF_X1 R2_temp_mix_data_reg_77_ ( .D(R2_n464), .CK(clk), .Q(R2_n302) );
  DLH_X1 R2_add_in_data_reg_76_ ( .G(R2_n2404), .D(R2_n301), .Q(R2_n948) );
  DFF_X1 R2_temp_mix_data_reg_76_ ( .D(R2_n463), .CK(clk), .Q(R2_n301) );
  DLH_X1 R2_add_in_data_reg_75_ ( .G(R2_n2398), .D(R2_n300), .Q(R2_n947) );
  DFF_X1 R2_temp_mix_data_reg_75_ ( .D(R2_n462), .CK(clk), .Q(R2_n300) );
  DLH_X1 R2_add_in_data_reg_74_ ( .G(R2_n2400), .D(R2_n299), .Q(R2_n946) );
  DFF_X1 R2_temp_mix_data_reg_74_ ( .D(R2_n461), .CK(clk), .Q(R2_n299) );
  DLH_X1 R2_add_in_data_reg_73_ ( .G(R2_n2399), .D(R2_n298), .Q(R2_n945) );
  DFF_X1 R2_temp_mix_data_reg_73_ ( .D(R2_n460), .CK(clk), .Q(R2_n298) );
  DLH_X1 R2_add_in_data_reg_72_ ( .G(R2_U23_Z_1), .D(R2_n297), .Q(R2_n944) );
  DFF_X1 R2_temp_mix_data_reg_72_ ( .D(R2_n459), .CK(clk), .Q(R2_n297) );
  DLH_X1 R2_add_in_data_reg_71_ ( .G(R2_U23_Z_1), .D(R2_n296), .Q(R2_n943) );
  DFF_X1 R2_temp_mix_data_reg_71_ ( .D(R2_n458), .CK(clk), .Q(R2_n296) );
  DLH_X1 R2_add_in_data_reg_70_ ( .G(R2_n2398), .D(R2_n295), .Q(R2_n942) );
  DFF_X1 R2_temp_mix_data_reg_70_ ( .D(R2_n457), .CK(clk), .Q(R2_n295) );
  DLH_X1 R2_add_in_data_reg_69_ ( .G(R2_U23_Z_1), .D(R2_n294), .Q(R2_n941) );
  DFF_X1 R2_temp_mix_data_reg_69_ ( .D(R2_n456), .CK(clk), .Q(R2_n294) );
  DLH_X1 R2_add_in_data_reg_68_ ( .G(R2_n2398), .D(R2_n293), .Q(R2_n940) );
  DFF_X1 R2_temp_mix_data_reg_68_ ( .D(R2_n455), .CK(clk), .Q(R2_n293) );
  DLH_X1 R2_add_in_data_reg_67_ ( .G(R2_n2403), .D(R2_n292), .Q(R2_n939) );
  DFF_X1 R2_temp_mix_data_reg_67_ ( .D(R2_n454), .CK(clk), .Q(R2_n292) );
  DLH_X1 R2_add_in_data_reg_66_ ( .G(R2_U23_Z_1), .D(R2_n291), .Q(R2_n938) );
  DFF_X1 R2_temp_mix_data_reg_66_ ( .D(R2_n453), .CK(clk), .Q(R2_n291) );
  DLH_X1 R2_add_in_data_reg_65_ ( .G(R2_n2401), .D(R2_n290), .Q(R2_n937) );
  DFF_X1 R2_temp_mix_data_reg_65_ ( .D(R2_n452), .CK(clk), .Q(R2_n290) );
  DLH_X1 R2_add_in_data_reg_64_ ( .G(R2_n2402), .D(R2_n289), .Q(R2_n936) );
  DFF_X1 R2_temp_mix_data_reg_64_ ( .D(R2_n451), .CK(clk), .Q(R2_n289) );
  DLH_X1 R2_add_in_data_reg_63_ ( .G(R2_n2402), .D(R2_n288), .Q(R2_n935) );
  DFF_X1 R2_temp_mix_data_reg_63_ ( .D(R2_n450), .CK(clk), .Q(R2_n288) );
  DLH_X1 R2_add_in_data_reg_62_ ( .G(R2_U23_Z_1), .D(R2_n287), .Q(R2_n934) );
  DFF_X1 R2_temp_mix_data_reg_62_ ( .D(R2_n449), .CK(clk), .Q(R2_n287) );
  DLH_X1 R2_add_in_data_reg_61_ ( .G(R2_n2402), .D(R2_n286), .Q(R2_n933) );
  DFF_X1 R2_temp_mix_data_reg_61_ ( .D(R2_n448), .CK(clk), .Q(R2_n286) );
  DLH_X1 R2_add_in_data_reg_60_ ( .G(R2_n2399), .D(R2_n285), .Q(R2_n932) );
  DFF_X1 R2_temp_mix_data_reg_60_ ( .D(R2_n447), .CK(clk), .Q(R2_n285) );
  DLH_X1 R2_add_in_data_reg_59_ ( .G(R2_n2398), .D(R2_n284), .Q(R2_n931) );
  DFF_X1 R2_temp_mix_data_reg_59_ ( .D(R2_n446), .CK(clk), .Q(R2_n284) );
  DLH_X1 R2_add_in_data_reg_58_ ( .G(R2_n2399), .D(R2_n283), .Q(R2_n930) );
  DFF_X1 R2_temp_mix_data_reg_58_ ( .D(R2_n445), .CK(clk), .Q(R2_n283) );
  DLH_X1 R2_add_in_data_reg_57_ ( .G(R2_U23_Z_1), .D(R2_n282), .Q(R2_n929) );
  DFF_X1 R2_temp_mix_data_reg_57_ ( .D(R2_n444), .CK(clk), .Q(R2_n282) );
  DLH_X1 R2_add_in_data_reg_56_ ( .G(R2_n2399), .D(R2_n281), .Q(R2_n928) );
  DFF_X1 R2_temp_mix_data_reg_56_ ( .D(R2_n443), .CK(clk), .Q(R2_n281) );
  DLH_X1 R2_add_in_data_reg_55_ ( .G(R2_n2401), .D(R2_n280), .Q(R2_n927) );
  DFF_X1 R2_temp_mix_data_reg_55_ ( .D(R2_n442), .CK(clk), .Q(R2_n280) );
  DLH_X1 R2_add_in_data_reg_54_ ( .G(R2_n2399), .D(R2_n279), .Q(R2_n926) );
  DFF_X1 R2_temp_mix_data_reg_54_ ( .D(R2_n441), .CK(clk), .Q(R2_n279) );
  DLH_X1 R2_add_in_data_reg_53_ ( .G(R2_n2402), .D(R2_n278), .Q(R2_n925) );
  DFF_X1 R2_temp_mix_data_reg_53_ ( .D(R2_n440), .CK(clk), .Q(R2_n278) );
  DLH_X1 R2_add_in_data_reg_52_ ( .G(R2_n2404), .D(R2_n277), .Q(R2_n924) );
  DFF_X1 R2_temp_mix_data_reg_52_ ( .D(R2_n439), .CK(clk), .Q(R2_n277) );
  DLH_X1 R2_add_in_data_reg_51_ ( .G(R2_n2402), .D(R2_n276), .Q(R2_n923) );
  DFF_X1 R2_temp_mix_data_reg_51_ ( .D(R2_n438), .CK(clk), .Q(R2_n276) );
  DLH_X1 R2_add_in_data_reg_50_ ( .G(R2_n2402), .D(R2_n275), .Q(R2_n922) );
  DFF_X1 R2_temp_mix_data_reg_50_ ( .D(R2_n437), .CK(clk), .Q(R2_n275) );
  DLH_X1 R2_add_in_data_reg_49_ ( .G(R2_n2403), .D(R2_n274), .Q(R2_n921) );
  DFF_X1 R2_temp_mix_data_reg_49_ ( .D(R2_n436), .CK(clk), .Q(R2_n274) );
  DLH_X1 R2_add_in_data_reg_48_ ( .G(R2_n2398), .D(R2_n273), .Q(R2_n920) );
  DFF_X1 R2_temp_mix_data_reg_48_ ( .D(R2_n435), .CK(clk), .Q(R2_n273) );
  DLH_X1 R2_add_in_data_reg_47_ ( .G(R2_n2403), .D(R2_n272), .Q(R2_n919) );
  DFF_X1 R2_temp_mix_data_reg_47_ ( .D(R2_n434), .CK(clk), .Q(R2_n272) );
  DLH_X1 R2_add_in_data_reg_46_ ( .G(R2_n2400), .D(R2_n271), .Q(R2_n918) );
  DFF_X1 R2_temp_mix_data_reg_46_ ( .D(R2_n433), .CK(clk), .Q(R2_n271) );
  DLH_X1 R2_add_in_data_reg_45_ ( .G(R2_n2398), .D(R2_n270), .Q(R2_n917) );
  DFF_X1 R2_temp_mix_data_reg_45_ ( .D(R2_n432), .CK(clk), .Q(R2_n270) );
  DLH_X1 R2_add_in_data_reg_44_ ( .G(R2_n2400), .D(R2_n269), .Q(R2_n916) );
  DFF_X1 R2_temp_mix_data_reg_44_ ( .D(R2_n431), .CK(clk), .Q(R2_n269) );
  DLH_X1 R2_add_in_data_reg_43_ ( .G(R2_n2404), .D(R2_n268), .Q(R2_n915) );
  DFF_X1 R2_temp_mix_data_reg_43_ ( .D(R2_n430), .CK(clk), .Q(R2_n268) );
  DLH_X1 R2_add_in_data_reg_42_ ( .G(R2_n2403), .D(R2_n267), .Q(R2_n914) );
  DFF_X1 R2_temp_mix_data_reg_42_ ( .D(R2_n429), .CK(clk), .Q(R2_n267) );
  DLH_X1 R2_add_in_data_reg_41_ ( .G(R2_n2400), .D(R2_n266), .Q(R2_n913) );
  DFF_X1 R2_temp_mix_data_reg_41_ ( .D(R2_n428), .CK(clk), .Q(R2_n266) );
  DLH_X1 R2_add_in_data_reg_40_ ( .G(R2_n2400), .D(R2_n265), .Q(R2_n912) );
  DFF_X1 R2_temp_mix_data_reg_40_ ( .D(R2_n427), .CK(clk), .Q(R2_n265) );
  DLH_X1 R2_add_in_data_reg_39_ ( .G(R2_n2402), .D(R2_n264), .Q(R2_n911) );
  DFF_X1 R2_temp_mix_data_reg_39_ ( .D(R2_n426), .CK(clk), .Q(R2_n264) );
  DLH_X1 R2_add_in_data_reg_38_ ( .G(R2_n2401), .D(R2_n263), .Q(R2_n910) );
  DFF_X1 R2_temp_mix_data_reg_38_ ( .D(R2_n425), .CK(clk), .Q(R2_n263) );
  DLH_X1 R2_add_in_data_reg_37_ ( .G(R2_n2401), .D(R2_n262), .Q(R2_n909) );
  DFF_X1 R2_temp_mix_data_reg_37_ ( .D(R2_n424), .CK(clk), .Q(R2_n262) );
  DLH_X1 R2_add_in_data_reg_36_ ( .G(R2_n2404), .D(R2_n261), .Q(R2_n908) );
  DFF_X1 R2_temp_mix_data_reg_36_ ( .D(R2_n423), .CK(clk), .Q(R2_n261) );
  DLH_X1 R2_add_in_data_reg_35_ ( .G(R2_n2404), .D(R2_n260), .Q(R2_n907) );
  DFF_X1 R2_temp_mix_data_reg_35_ ( .D(R2_n422), .CK(clk), .Q(R2_n260) );
  DLH_X1 R2_add_in_data_reg_34_ ( .G(R2_U23_Z_1), .D(R2_n259), .Q(R2_n906) );
  DFF_X1 R2_temp_mix_data_reg_34_ ( .D(R2_n421), .CK(clk), .Q(R2_n259) );
  DLH_X1 R2_add_in_data_reg_33_ ( .G(R2_n2402), .D(R2_n258), .Q(R2_n905) );
  DFF_X1 R2_temp_mix_data_reg_33_ ( .D(R2_n420), .CK(clk), .Q(R2_n258) );
  DLH_X1 R2_add_in_data_reg_32_ ( .G(R2_n2403), .D(R2_n257), .Q(R2_n904) );
  DFF_X1 R2_temp_mix_data_reg_32_ ( .D(R2_n419), .CK(clk), .Q(R2_n257) );
  DLH_X1 R2_add_in_data_reg_31_ ( .G(R2_n2401), .D(R2_n256), .Q(R2_n903) );
  DFF_X1 R2_temp_mix_data_reg_31_ ( .D(R2_n418), .CK(clk), .Q(R2_n256) );
  DLH_X1 R2_add_in_data_reg_30_ ( .G(R2_n2399), .D(R2_n255), .Q(R2_n902) );
  DFF_X1 R2_temp_mix_data_reg_30_ ( .D(R2_n417), .CK(clk), .Q(R2_n255) );
  DLH_X1 R2_add_in_data_reg_29_ ( .G(R2_n2401), .D(R2_n254), .Q(R2_n901) );
  DFF_X1 R2_temp_mix_data_reg_29_ ( .D(R2_n416), .CK(clk), .Q(R2_n254) );
  DLH_X1 R2_add_in_data_reg_28_ ( .G(R2_n2399), .D(R2_n253), .Q(R2_n900) );
  DFF_X1 R2_temp_mix_data_reg_28_ ( .D(R2_n415), .CK(clk), .Q(R2_n253) );
  DLH_X1 R2_add_in_data_reg_27_ ( .G(R2_U23_Z_1), .D(R2_n252), .Q(R2_n899) );
  DFF_X1 R2_temp_mix_data_reg_27_ ( .D(R2_n414), .CK(clk), .Q(R2_n252) );
  DLH_X1 R2_add_in_data_reg_26_ ( .G(R2_n2400), .D(R2_n251), .Q(R2_n898) );
  DFF_X1 R2_temp_mix_data_reg_26_ ( .D(R2_n413), .CK(clk), .Q(R2_n251) );
  DLH_X1 R2_add_in_data_reg_25_ ( .G(R2_U23_Z_1), .D(R2_n250), .Q(R2_n897) );
  DFF_X1 R2_temp_mix_data_reg_25_ ( .D(R2_n412), .CK(clk), .Q(R2_n250) );
  DLH_X1 R2_add_in_data_reg_24_ ( .G(R2_n2398), .D(R2_n249), .Q(R2_n896) );
  DFF_X1 R2_temp_mix_data_reg_24_ ( .D(R2_n411), .CK(clk), .Q(R2_n249) );
  DLH_X1 R2_add_in_data_reg_23_ ( .G(R2_U23_Z_1), .D(R2_n248), .Q(R2_n895) );
  DFF_X1 R2_temp_mix_data_reg_23_ ( .D(R2_n410), .CK(clk), .Q(R2_n248) );
  DLH_X1 R2_add_in_data_reg_22_ ( .G(R2_n2398), .D(R2_n247), .Q(R2_n894) );
  DFF_X1 R2_temp_mix_data_reg_22_ ( .D(R2_n409), .CK(clk), .Q(R2_n247) );
  DLH_X1 R2_add_in_data_reg_21_ ( .G(R2_n2398), .D(R2_n246), .Q(R2_n893) );
  DFF_X1 R2_temp_mix_data_reg_21_ ( .D(R2_n408), .CK(clk), .Q(R2_n246) );
  DLH_X1 R2_add_in_data_reg_20_ ( .G(R2_n2402), .D(R2_n245), .Q(R2_n892) );
  DFF_X1 R2_temp_mix_data_reg_20_ ( .D(R2_n407), .CK(clk), .Q(R2_n245) );
  DLH_X1 R2_add_in_data_reg_19_ ( .G(R2_U23_Z_1), .D(R2_n244), .Q(R2_n891) );
  DFF_X1 R2_temp_mix_data_reg_19_ ( .D(R2_n406), .CK(clk), .Q(R2_n244) );
  DLH_X1 R2_add_in_data_reg_18_ ( .G(R2_n2400), .D(R2_n243), .Q(R2_n890) );
  DFF_X1 R2_temp_mix_data_reg_18_ ( .D(R2_n405), .CK(clk), .Q(R2_n243) );
  DLH_X1 R2_add_in_data_reg_17_ ( .G(R2_n2401), .D(R2_n242), .Q(R2_n889) );
  DFF_X1 R2_temp_mix_data_reg_17_ ( .D(R2_n404), .CK(clk), .Q(R2_n242) );
  DLH_X1 R2_add_in_data_reg_16_ ( .G(R2_n2403), .D(R2_n241), .Q(R2_n888) );
  DFF_X1 R2_temp_mix_data_reg_16_ ( .D(R2_n403), .CK(clk), .Q(R2_n241) );
  DLH_X1 R2_add_in_data_reg_15_ ( .G(R2_n2400), .D(R2_n240), .Q(R2_n887) );
  DFF_X1 R2_temp_mix_data_reg_15_ ( .D(R2_n402), .CK(clk), .Q(R2_n240) );
  DLH_X1 R2_add_in_data_reg_14_ ( .G(R2_n2403), .D(R2_n239), .Q(R2_n886) );
  DFF_X1 R2_temp_mix_data_reg_14_ ( .D(R2_n401), .CK(clk), .Q(R2_n239) );
  DLH_X1 R2_add_in_data_reg_13_ ( .G(R2_n2400), .D(R2_n238), .Q(R2_n885) );
  DFF_X1 R2_temp_mix_data_reg_13_ ( .D(R2_n400), .CK(clk), .Q(R2_n238) );
  DLH_X1 R2_add_in_data_reg_12_ ( .G(R2_n2401), .D(R2_n237), .Q(R2_n884) );
  DFF_X1 R2_temp_mix_data_reg_12_ ( .D(R2_n399), .CK(clk), .Q(R2_n237) );
  DLH_X1 R2_add_in_data_reg_11_ ( .G(R2_n2403), .D(R2_n236), .Q(R2_n883) );
  DFF_X1 R2_temp_mix_data_reg_11_ ( .D(R2_n398), .CK(clk), .Q(R2_n236) );
  DLH_X1 R2_add_in_data_reg_10_ ( .G(R2_n2402), .D(R2_n235), .Q(R2_n882) );
  DFF_X1 R2_temp_mix_data_reg_10_ ( .D(R2_n397), .CK(clk), .Q(R2_n235) );
  DLH_X1 R2_add_in_data_reg_9_ ( .G(R2_n2399), .D(R2_n234), .Q(R2_n881) );
  DFF_X1 R2_temp_mix_data_reg_9_ ( .D(R2_n396), .CK(clk), .Q(R2_n234) );
  DLH_X1 R2_add_in_data_reg_8_ ( .G(R2_n2404), .D(R2_n233), .Q(R2_n880) );
  DFF_X1 R2_temp_mix_data_reg_8_ ( .D(R2_n395), .CK(clk), .Q(R2_n233) );
  DLH_X1 R2_add_in_data_reg_7_ ( .G(R2_n2401), .D(R2_n232), .Q(R2_n879) );
  DFF_X1 R2_temp_mix_data_reg_7_ ( .D(R2_n394), .CK(clk), .Q(R2_n232) );
  DLH_X1 R2_add_in_data_reg_6_ ( .G(R2_n2403), .D(R2_n231), .Q(R2_n878) );
  DFF_X1 R2_temp_mix_data_reg_6_ ( .D(R2_n393), .CK(clk), .Q(R2_n231) );
  DLH_X1 R2_add_in_data_reg_5_ ( .G(R2_n2400), .D(R2_n230), .Q(R2_n877) );
  DFF_X1 R2_temp_mix_data_reg_5_ ( .D(R2_n392), .CK(clk), .Q(R2_n230) );
  DLH_X1 R2_add_in_data_reg_4_ ( .G(R2_n2404), .D(R2_n229), .Q(R2_n876) );
  DFF_X1 R2_temp_mix_data_reg_4_ ( .D(R2_n391), .CK(clk), .Q(R2_n229) );
  DLH_X1 R2_add_in_data_reg_3_ ( .G(R2_n2401), .D(R2_n228), .Q(R2_n875) );
  DFF_X1 R2_temp_mix_data_reg_3_ ( .D(R2_n390), .CK(clk), .Q(R2_n228) );
  DLH_X1 R2_add_in_data_reg_2_ ( .G(R2_U23_Z_1), .D(R2_n227), .Q(R2_n874) );
  DFF_X1 R2_temp_mix_data_reg_2_ ( .D(R2_n389), .CK(clk), .Q(R2_n227) );
  DLH_X1 R2_add_in_data_reg_1_ ( .G(R2_n2398), .D(R2_n226), .Q(R2_n873) );
  DFF_X1 R2_temp_mix_data_reg_1_ ( .D(R2_n388), .CK(clk), .Q(R2_n226) );
  DLH_X1 R2_add_in_data_reg_0_ ( .G(R2_n2404), .D(R2_n225), .Q(R2_n872) );
  DFF_X1 R2_temp_mix_data_reg_0_ ( .D(R2_n387), .CK(clk), .Q(R2_n225) );
  DLH_X1 R2_mix_in_data_reg_127_ ( .G(R2_n2394), .D(R2_U16_DATA1_127), .Q(
        R2_n1256) );
  DFF_X1 R2_temp_shift_data_reg_127_ ( .D(R2_n386), .CK(clk), .Q(
        R2_U16_DATA1_127) );
  DLH_X1 R2_mix_in_data_reg_126_ ( .G(R2_n2394), .D(R2_U16_DATA1_126), .Q(
        R2_n1255) );
  DFF_X1 R2_temp_shift_data_reg_126_ ( .D(R2_n385), .CK(clk), .Q(
        R2_U16_DATA1_126) );
  DLH_X1 R2_mix_in_data_reg_125_ ( .G(R2_n2392), .D(R2_U16_DATA1_125), .Q(
        R2_n1254) );
  DFF_X1 R2_temp_shift_data_reg_125_ ( .D(R2_n384), .CK(clk), .Q(
        R2_U16_DATA1_125) );
  DLH_X1 R2_mix_in_data_reg_124_ ( .G(R2_n2393), .D(R2_U16_DATA1_124), .Q(
        R2_n1253) );
  DFF_X1 R2_temp_shift_data_reg_124_ ( .D(R2_n383), .CK(clk), .Q(
        R2_U16_DATA1_124) );
  DLH_X1 R2_mix_in_data_reg_123_ ( .G(R2_n2391), .D(R2_U16_DATA1_123), .Q(
        R2_n1252) );
  DFF_X1 R2_temp_shift_data_reg_123_ ( .D(R2_n382), .CK(clk), .Q(
        R2_U16_DATA1_123) );
  DLH_X1 R2_mix_in_data_reg_122_ ( .G(R2_n2391), .D(R2_U16_DATA1_122), .Q(
        R2_n1251) );
  DFF_X1 R2_temp_shift_data_reg_122_ ( .D(R2_n381), .CK(clk), .Q(
        R2_U16_DATA1_122) );
  DLH_X1 R2_mix_in_data_reg_121_ ( .G(R2_n2393), .D(R2_U16_DATA1_121), .Q(
        R2_n1250) );
  DFF_X1 R2_temp_shift_data_reg_121_ ( .D(R2_n380), .CK(clk), .Q(
        R2_U16_DATA1_121) );
  DLH_X1 R2_mix_in_data_reg_120_ ( .G(R2_n2394), .D(R2_U16_DATA1_120), .Q(
        R2_n1249) );
  DFF_X1 R2_temp_shift_data_reg_120_ ( .D(R2_n379), .CK(clk), .Q(
        R2_U16_DATA1_120) );
  DLH_X1 R2_mix_in_data_reg_119_ ( .G(R2_n2391), .D(R2_U16_DATA1_119), .Q(
        R2_n1248) );
  DFF_X1 R2_temp_shift_data_reg_119_ ( .D(R2_n378), .CK(clk), .Q(
        R2_U16_DATA1_119) );
  DLH_X1 R2_mix_in_data_reg_118_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_118), .Q(
        R2_n1247) );
  DFF_X1 R2_temp_shift_data_reg_118_ ( .D(R2_n377), .CK(clk), .Q(
        R2_U16_DATA1_118) );
  DLH_X1 R2_mix_in_data_reg_117_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_117), .Q(
        R2_n1246) );
  DFF_X1 R2_temp_shift_data_reg_117_ ( .D(R2_n376), .CK(clk), .Q(
        R2_U16_DATA1_117) );
  DLH_X1 R2_mix_in_data_reg_116_ ( .G(R2_n2394), .D(R2_U16_DATA1_116), .Q(
        R2_n1245) );
  DFF_X1 R2_temp_shift_data_reg_116_ ( .D(R2_n375), .CK(clk), .Q(
        R2_U16_DATA1_116) );
  DLH_X1 R2_mix_in_data_reg_115_ ( .G(R2_n2392), .D(R2_U16_DATA1_115), .Q(
        R2_n1244) );
  DFF_X1 R2_temp_shift_data_reg_115_ ( .D(R2_n374), .CK(clk), .Q(
        R2_U16_DATA1_115) );
  DLH_X1 R2_mix_in_data_reg_114_ ( .G(R2_n2391), .D(R2_U16_DATA1_114), .Q(
        R2_n1243) );
  DFF_X1 R2_temp_shift_data_reg_114_ ( .D(R2_n373), .CK(clk), .Q(
        R2_U16_DATA1_114) );
  DLH_X1 R2_mix_in_data_reg_113_ ( .G(R2_n2394), .D(R2_U16_DATA1_113), .Q(
        R2_n1242) );
  DFF_X1 R2_temp_shift_data_reg_113_ ( .D(R2_n372), .CK(clk), .Q(
        R2_U16_DATA1_113) );
  DLH_X1 R2_mix_in_data_reg_112_ ( .G(R2_n2394), .D(R2_U16_DATA1_112), .Q(
        R2_n1241) );
  DFF_X1 R2_temp_shift_data_reg_112_ ( .D(R2_n371), .CK(clk), .Q(
        R2_U16_DATA1_112) );
  DLH_X1 R2_mix_in_data_reg_111_ ( .G(R2_n2393), .D(R2_U16_DATA1_111), .Q(
        R2_n1240) );
  DFF_X1 R2_temp_shift_data_reg_111_ ( .D(R2_n370), .CK(clk), .Q(
        R2_U16_DATA1_111) );
  DLH_X1 R2_mix_in_data_reg_110_ ( .G(R2_n2392), .D(R2_U16_DATA1_110), .Q(
        R2_n1239) );
  DFF_X1 R2_temp_shift_data_reg_110_ ( .D(R2_n369), .CK(clk), .Q(
        R2_U16_DATA1_110) );
  DLH_X1 R2_mix_in_data_reg_109_ ( .G(R2_n2394), .D(R2_U16_DATA1_109), .Q(
        R2_n1238) );
  DFF_X1 R2_temp_shift_data_reg_109_ ( .D(R2_n368), .CK(clk), .Q(
        R2_U16_DATA1_109) );
  DLH_X1 R2_mix_in_data_reg_108_ ( .G(R2_n2391), .D(R2_U16_DATA1_108), .Q(
        R2_n1237) );
  DFF_X1 R2_temp_shift_data_reg_108_ ( .D(R2_n367), .CK(clk), .Q(
        R2_U16_DATA1_108) );
  DLH_X1 R2_mix_in_data_reg_107_ ( .G(R2_n2392), .D(R2_U16_DATA1_107), .Q(
        R2_n1236) );
  DFF_X1 R2_temp_shift_data_reg_107_ ( .D(R2_n366), .CK(clk), .Q(
        R2_U16_DATA1_107) );
  DLH_X1 R2_mix_in_data_reg_106_ ( .G(R2_n2393), .D(R2_U16_DATA1_106), .Q(
        R2_n1235) );
  DFF_X1 R2_temp_shift_data_reg_106_ ( .D(R2_n365), .CK(clk), .Q(
        R2_U16_DATA1_106) );
  DLH_X1 R2_mix_in_data_reg_105_ ( .G(R2_n2392), .D(R2_U16_DATA1_105), .Q(
        R2_n1234) );
  DFF_X1 R2_temp_shift_data_reg_105_ ( .D(R2_n364), .CK(clk), .Q(
        R2_U16_DATA1_105) );
  DLH_X1 R2_mix_in_data_reg_104_ ( .G(R2_n2392), .D(R2_U16_DATA1_104), .Q(
        R2_n1233) );
  DFF_X1 R2_temp_shift_data_reg_104_ ( .D(R2_n363), .CK(clk), .Q(
        R2_U16_DATA1_104) );
  DLH_X1 R2_mix_in_data_reg_103_ ( .G(R2_n2393), .D(R2_U16_DATA1_103), .Q(
        R2_n1232) );
  DFF_X1 R2_temp_shift_data_reg_103_ ( .D(R2_n362), .CK(clk), .Q(
        R2_U16_DATA1_103) );
  DLH_X1 R2_mix_in_data_reg_102_ ( .G(R2_n2393), .D(R2_U16_DATA1_102), .Q(
        R2_n1231) );
  DFF_X1 R2_temp_shift_data_reg_102_ ( .D(R2_n361), .CK(clk), .Q(
        R2_U16_DATA1_102) );
  DLH_X1 R2_mix_in_data_reg_101_ ( .G(R2_n2394), .D(R2_U16_DATA1_101), .Q(
        R2_n1230) );
  DFF_X1 R2_temp_shift_data_reg_101_ ( .D(R2_n360), .CK(clk), .Q(
        R2_U16_DATA1_101) );
  DLH_X1 R2_mix_in_data_reg_100_ ( .G(R2_n2393), .D(R2_U16_DATA1_100), .Q(
        R2_n1229) );
  DFF_X1 R2_temp_shift_data_reg_100_ ( .D(R2_n359), .CK(clk), .Q(
        R2_U16_DATA1_100) );
  DLH_X1 R2_mix_in_data_reg_99_ ( .G(R2_n2394), .D(R2_U16_DATA1_99), .Q(
        R2_n1228) );
  DFF_X1 R2_temp_shift_data_reg_99_ ( .D(R2_n358), .CK(clk), .Q(
        R2_U16_DATA1_99) );
  DLH_X1 R2_mix_in_data_reg_98_ ( .G(R2_n2391), .D(R2_U16_DATA1_98), .Q(
        R2_n1227) );
  DFF_X1 R2_temp_shift_data_reg_98_ ( .D(R2_n357), .CK(clk), .Q(
        R2_U16_DATA1_98) );
  DLH_X1 R2_mix_in_data_reg_97_ ( .G(R2_n2391), .D(R2_U16_DATA1_97), .Q(
        R2_n1226) );
  DFF_X1 R2_temp_shift_data_reg_97_ ( .D(R2_n356), .CK(clk), .Q(
        R2_U16_DATA1_97) );
  DLH_X1 R2_mix_in_data_reg_96_ ( .G(R2_n2391), .D(R2_U16_DATA1_96), .Q(
        R2_n1225) );
  DFF_X1 R2_temp_shift_data_reg_96_ ( .D(R2_n355), .CK(clk), .Q(
        R2_U16_DATA1_96) );
  DLH_X1 R2_mix_in_data_reg_95_ ( .G(R2_n2393), .D(R2_U16_DATA1_95), .Q(
        R2_n1224) );
  DFF_X1 R2_temp_shift_data_reg_95_ ( .D(R2_n354), .CK(clk), .Q(
        R2_U16_DATA1_95) );
  DLH_X1 R2_mix_in_data_reg_94_ ( .G(R2_n2393), .D(R2_U16_DATA1_94), .Q(
        R2_n1223) );
  DFF_X1 R2_temp_shift_data_reg_94_ ( .D(R2_n353), .CK(clk), .Q(
        R2_U16_DATA1_94) );
  DLH_X1 R2_mix_in_data_reg_93_ ( .G(R2_n2391), .D(R2_U16_DATA1_93), .Q(
        R2_n1222) );
  DFF_X1 R2_temp_shift_data_reg_93_ ( .D(R2_n224), .CK(clk), .Q(
        R2_U16_DATA1_93) );
  DLH_X1 R2_mix_in_data_reg_92_ ( .G(R2_n2392), .D(R2_U16_DATA1_92), .Q(
        R2_n1221) );
  DFF_X1 R2_temp_shift_data_reg_92_ ( .D(R2_n223), .CK(clk), .Q(
        R2_U16_DATA1_92) );
  DLH_X1 R2_mix_in_data_reg_91_ ( .G(R2_n2391), .D(R2_U16_DATA1_91), .Q(
        R2_n1220) );
  DFF_X1 R2_temp_shift_data_reg_91_ ( .D(R2_n222), .CK(clk), .Q(
        R2_U16_DATA1_91) );
  DLH_X1 R2_mix_in_data_reg_90_ ( .G(R2_n2393), .D(R2_U16_DATA1_90), .Q(
        R2_n1219) );
  DFF_X1 R2_temp_shift_data_reg_90_ ( .D(R2_n221), .CK(clk), .Q(
        R2_U16_DATA1_90) );
  DLH_X1 R2_mix_in_data_reg_89_ ( .G(R2_n2391), .D(R2_U16_DATA1_89), .Q(
        R2_n1218) );
  DFF_X1 R2_temp_shift_data_reg_89_ ( .D(R2_n220), .CK(clk), .Q(
        R2_U16_DATA1_89) );
  DLH_X1 R2_mix_in_data_reg_88_ ( .G(R2_n2392), .D(R2_U16_DATA1_88), .Q(
        R2_n1217) );
  DFF_X1 R2_temp_shift_data_reg_88_ ( .D(R2_n219), .CK(clk), .Q(
        R2_U16_DATA1_88) );
  DLH_X1 R2_mix_in_data_reg_87_ ( .G(R2_n2394), .D(R2_U16_DATA1_87), .Q(
        R2_n1216) );
  DFF_X1 R2_temp_shift_data_reg_87_ ( .D(R2_n218), .CK(clk), .Q(
        R2_U16_DATA1_87) );
  DLH_X1 R2_mix_in_data_reg_86_ ( .G(R2_n2393), .D(R2_U16_DATA1_86), .Q(
        R2_n1215) );
  DFF_X1 R2_temp_shift_data_reg_86_ ( .D(R2_n217), .CK(clk), .Q(
        R2_U16_DATA1_86) );
  DLH_X1 R2_mix_in_data_reg_85_ ( .G(R2_n2394), .D(R2_U16_DATA1_85), .Q(
        R2_n1214) );
  DFF_X1 R2_temp_shift_data_reg_85_ ( .D(R2_n216), .CK(clk), .Q(
        R2_U16_DATA1_85) );
  DLH_X1 R2_mix_in_data_reg_84_ ( .G(R2_n2393), .D(R2_U16_DATA1_84), .Q(
        R2_n1213) );
  DFF_X1 R2_temp_shift_data_reg_84_ ( .D(R2_n215), .CK(clk), .Q(
        R2_U16_DATA1_84) );
  DLH_X1 R2_mix_in_data_reg_83_ ( .G(R2_n2392), .D(R2_U16_DATA1_83), .Q(
        R2_n1212) );
  DFF_X1 R2_temp_shift_data_reg_83_ ( .D(R2_n214), .CK(clk), .Q(
        R2_U16_DATA1_83) );
  DLH_X1 R2_mix_in_data_reg_82_ ( .G(R2_n2393), .D(R2_U16_DATA1_82), .Q(
        R2_n1211) );
  DFF_X1 R2_temp_shift_data_reg_82_ ( .D(R2_n213), .CK(clk), .Q(
        R2_U16_DATA1_82) );
  DLH_X1 R2_mix_in_data_reg_81_ ( .G(R2_n2393), .D(R2_U16_DATA1_81), .Q(
        R2_n1210) );
  DFF_X1 R2_temp_shift_data_reg_81_ ( .D(R2_n212), .CK(clk), .Q(
        R2_U16_DATA1_81) );
  DLH_X1 R2_mix_in_data_reg_80_ ( .G(R2_n2391), .D(R2_U16_DATA1_80), .Q(
        R2_n1209) );
  DFF_X1 R2_temp_shift_data_reg_80_ ( .D(R2_n211), .CK(clk), .Q(
        R2_U16_DATA1_80) );
  DLH_X1 R2_mix_in_data_reg_79_ ( .G(R2_n2394), .D(R2_U16_DATA1_79), .Q(
        R2_n1208) );
  DFF_X1 R2_temp_shift_data_reg_79_ ( .D(R2_n210), .CK(clk), .Q(
        R2_U16_DATA1_79) );
  DLH_X1 R2_mix_in_data_reg_78_ ( .G(R2_n2391), .D(R2_U16_DATA1_78), .Q(
        R2_n1207) );
  DFF_X1 R2_temp_shift_data_reg_78_ ( .D(R2_n209), .CK(clk), .Q(
        R2_U16_DATA1_78) );
  DLH_X1 R2_mix_in_data_reg_77_ ( .G(R2_n2392), .D(R2_U16_DATA1_77), .Q(
        R2_n1206) );
  DFF_X1 R2_temp_shift_data_reg_77_ ( .D(R2_n208), .CK(clk), .Q(
        R2_U16_DATA1_77) );
  DLH_X1 R2_mix_in_data_reg_76_ ( .G(R2_n2391), .D(R2_U16_DATA1_76), .Q(
        R2_n1205) );
  DFF_X1 R2_temp_shift_data_reg_76_ ( .D(R2_n207), .CK(clk), .Q(
        R2_U16_DATA1_76) );
  DLH_X1 R2_mix_in_data_reg_75_ ( .G(R2_n2393), .D(R2_U16_DATA1_75), .Q(
        R2_n1204) );
  DFF_X1 R2_temp_shift_data_reg_75_ ( .D(R2_n206), .CK(clk), .Q(
        R2_U16_DATA1_75) );
  DLH_X1 R2_mix_in_data_reg_74_ ( .G(R2_n2392), .D(R2_U16_DATA1_74), .Q(
        R2_n1203) );
  DFF_X1 R2_temp_shift_data_reg_74_ ( .D(R2_n205), .CK(clk), .Q(
        R2_U16_DATA1_74) );
  DLH_X1 R2_mix_in_data_reg_73_ ( .G(R2_n2394), .D(R2_U16_DATA1_73), .Q(
        R2_n1202) );
  DFF_X1 R2_temp_shift_data_reg_73_ ( .D(R2_n204), .CK(clk), .Q(
        R2_U16_DATA1_73) );
  DLH_X1 R2_mix_in_data_reg_72_ ( .G(R2_n2391), .D(R2_U16_DATA1_72), .Q(
        R2_n1201) );
  DFF_X1 R2_temp_shift_data_reg_72_ ( .D(R2_n203), .CK(clk), .Q(
        R2_U16_DATA1_72) );
  DLH_X1 R2_mix_in_data_reg_71_ ( .G(R2_n2392), .D(R2_U16_DATA1_71), .Q(
        R2_n1200) );
  DFF_X1 R2_temp_shift_data_reg_71_ ( .D(R2_n202), .CK(clk), .Q(
        R2_U16_DATA1_71) );
  DLH_X1 R2_mix_in_data_reg_70_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_70), .Q(
        R2_n1199) );
  DFF_X1 R2_temp_shift_data_reg_70_ ( .D(R2_n201), .CK(clk), .Q(
        R2_U16_DATA1_70) );
  DLH_X1 R2_mix_in_data_reg_69_ ( .G(R2_n2393), .D(R2_U16_DATA1_69), .Q(
        R2_n1198) );
  DFF_X1 R2_temp_shift_data_reg_69_ ( .D(R2_n200), .CK(clk), .Q(
        R2_U16_DATA1_69) );
  DLH_X1 R2_mix_in_data_reg_68_ ( .G(R2_n2392), .D(R2_U16_DATA1_68), .Q(
        R2_n1197) );
  DFF_X1 R2_temp_shift_data_reg_68_ ( .D(R2_n199), .CK(clk), .Q(
        R2_U16_DATA1_68) );
  DLH_X1 R2_mix_in_data_reg_67_ ( .G(R2_n2392), .D(R2_U16_DATA1_67), .Q(
        R2_n1196) );
  DFF_X1 R2_temp_shift_data_reg_67_ ( .D(R2_n198), .CK(clk), .Q(
        R2_U16_DATA1_67) );
  DLH_X1 R2_mix_in_data_reg_66_ ( .G(R2_n2393), .D(R2_U16_DATA1_66), .Q(
        R2_n1195) );
  DFF_X1 R2_temp_shift_data_reg_66_ ( .D(R2_n197), .CK(clk), .Q(
        R2_U16_DATA1_66) );
  DLH_X1 R2_mix_in_data_reg_65_ ( .G(R2_n2391), .D(R2_U16_DATA1_65), .Q(
        R2_n1194) );
  DFF_X1 R2_temp_shift_data_reg_65_ ( .D(R2_n196), .CK(clk), .Q(
        R2_U16_DATA1_65) );
  DLH_X1 R2_mix_in_data_reg_64_ ( .G(R2_n2394), .D(R2_U16_DATA1_64), .Q(
        R2_n1193) );
  DFF_X1 R2_temp_shift_data_reg_64_ ( .D(R2_n195), .CK(clk), .Q(
        R2_U16_DATA1_64) );
  DLH_X1 R2_mix_in_data_reg_63_ ( .G(R2_n2394), .D(R2_U16_DATA1_63), .Q(
        R2_n1192) );
  DFF_X1 R2_temp_shift_data_reg_63_ ( .D(R2_n194), .CK(clk), .Q(
        R2_U16_DATA1_63) );
  DLH_X1 R2_mix_in_data_reg_62_ ( .G(R2_n2391), .D(R2_U16_DATA1_62), .Q(
        R2_n1191) );
  DFF_X1 R2_temp_shift_data_reg_62_ ( .D(R2_n193), .CK(clk), .Q(
        R2_U16_DATA1_62) );
  DLH_X1 R2_mix_in_data_reg_61_ ( .G(R2_n2391), .D(R2_U16_DATA1_61), .Q(
        R2_n1190) );
  DFF_X1 R2_temp_shift_data_reg_61_ ( .D(R2_n192), .CK(clk), .Q(
        R2_U16_DATA1_61) );
  DLH_X1 R2_mix_in_data_reg_60_ ( .G(R2_n2391), .D(R2_U16_DATA1_60), .Q(
        R2_n1189) );
  DFF_X1 R2_temp_shift_data_reg_60_ ( .D(R2_n191), .CK(clk), .Q(
        R2_U16_DATA1_60) );
  DLH_X1 R2_mix_in_data_reg_59_ ( .G(R2_n2391), .D(R2_U16_DATA1_59), .Q(
        R2_n1188) );
  DFF_X1 R2_temp_shift_data_reg_59_ ( .D(R2_n190), .CK(clk), .Q(
        R2_U16_DATA1_59) );
  DLH_X1 R2_mix_in_data_reg_58_ ( .G(R2_n2391), .D(R2_U16_DATA1_58), .Q(
        R2_n1187) );
  DFF_X1 R2_temp_shift_data_reg_58_ ( .D(R2_n189), .CK(clk), .Q(
        R2_U16_DATA1_58) );
  DLH_X1 R2_mix_in_data_reg_57_ ( .G(R2_n2391), .D(R2_U16_DATA1_57), .Q(
        R2_n1186) );
  DFF_X1 R2_temp_shift_data_reg_57_ ( .D(R2_n188), .CK(clk), .Q(
        R2_U16_DATA1_57) );
  DLH_X1 R2_mix_in_data_reg_56_ ( .G(R2_n2391), .D(R2_U16_DATA1_56), .Q(
        R2_n1185) );
  DFF_X1 R2_temp_shift_data_reg_56_ ( .D(R2_n187), .CK(clk), .Q(
        R2_U16_DATA1_56) );
  DLH_X1 R2_mix_in_data_reg_55_ ( .G(R2_n2391), .D(R2_U16_DATA1_55), .Q(
        R2_n1184) );
  DFF_X1 R2_temp_shift_data_reg_55_ ( .D(R2_n186), .CK(clk), .Q(
        R2_U16_DATA1_55) );
  DLH_X1 R2_mix_in_data_reg_54_ ( .G(R2_n2391), .D(R2_U16_DATA1_54), .Q(
        R2_n1183) );
  DFF_X1 R2_temp_shift_data_reg_54_ ( .D(R2_n185), .CK(clk), .Q(
        R2_U16_DATA1_54) );
  DLH_X1 R2_mix_in_data_reg_53_ ( .G(R2_n2391), .D(R2_U16_DATA1_53), .Q(
        R2_n1182) );
  DFF_X1 R2_temp_shift_data_reg_53_ ( .D(R2_n184), .CK(clk), .Q(
        R2_U16_DATA1_53) );
  DLH_X1 R2_mix_in_data_reg_52_ ( .G(R2_n2391), .D(R2_U16_DATA1_52), .Q(
        R2_n1181) );
  DFF_X1 R2_temp_shift_data_reg_52_ ( .D(R2_n183), .CK(clk), .Q(
        R2_U16_DATA1_52) );
  DLH_X1 R2_mix_in_data_reg_51_ ( .G(R2_n2391), .D(R2_U16_DATA1_51), .Q(
        R2_n1180) );
  DFF_X1 R2_temp_shift_data_reg_51_ ( .D(R2_n182), .CK(clk), .Q(
        R2_U16_DATA1_51) );
  DLH_X1 R2_mix_in_data_reg_50_ ( .G(R2_n2392), .D(R2_U16_DATA1_50), .Q(
        R2_n1179) );
  DFF_X1 R2_temp_shift_data_reg_50_ ( .D(R2_n181), .CK(clk), .Q(
        R2_U16_DATA1_50) );
  DLH_X1 R2_mix_in_data_reg_49_ ( .G(R2_n2392), .D(R2_U16_DATA1_49), .Q(
        R2_n1178) );
  DFF_X1 R2_temp_shift_data_reg_49_ ( .D(R2_n180), .CK(clk), .Q(
        R2_U16_DATA1_49) );
  DLH_X1 R2_mix_in_data_reg_48_ ( .G(R2_n2392), .D(R2_U16_DATA1_48), .Q(
        R2_n1177) );
  DFF_X1 R2_temp_shift_data_reg_48_ ( .D(R2_n179), .CK(clk), .Q(
        R2_U16_DATA1_48) );
  DLH_X1 R2_mix_in_data_reg_47_ ( .G(R2_n2392), .D(R2_U16_DATA1_47), .Q(
        R2_n1176) );
  DFF_X1 R2_temp_shift_data_reg_47_ ( .D(R2_n178), .CK(clk), .Q(
        R2_U16_DATA1_47) );
  DLH_X1 R2_mix_in_data_reg_46_ ( .G(R2_n2392), .D(R2_U16_DATA1_46), .Q(
        R2_n1175) );
  DFF_X1 R2_temp_shift_data_reg_46_ ( .D(R2_n177), .CK(clk), .Q(
        R2_U16_DATA1_46) );
  DLH_X1 R2_mix_in_data_reg_45_ ( .G(R2_n2392), .D(R2_U16_DATA1_45), .Q(
        R2_n1174) );
  DFF_X1 R2_temp_shift_data_reg_45_ ( .D(R2_n176), .CK(clk), .Q(
        R2_U16_DATA1_45) );
  DLH_X1 R2_mix_in_data_reg_44_ ( .G(R2_n2392), .D(R2_U16_DATA1_44), .Q(
        R2_n1173) );
  DFF_X1 R2_temp_shift_data_reg_44_ ( .D(R2_n175), .CK(clk), .Q(
        R2_U16_DATA1_44) );
  DLH_X1 R2_mix_in_data_reg_43_ ( .G(R2_n2392), .D(R2_U16_DATA1_43), .Q(
        R2_n1172) );
  DFF_X1 R2_temp_shift_data_reg_43_ ( .D(R2_n174), .CK(clk), .Q(
        R2_U16_DATA1_43) );
  DLH_X1 R2_mix_in_data_reg_42_ ( .G(R2_n2392), .D(R2_U16_DATA1_42), .Q(
        R2_n1171) );
  DFF_X1 R2_temp_shift_data_reg_42_ ( .D(R2_n173), .CK(clk), .Q(
        R2_U16_DATA1_42) );
  DLH_X1 R2_mix_in_data_reg_41_ ( .G(R2_n2392), .D(R2_U16_DATA1_41), .Q(
        R2_n1170) );
  DFF_X1 R2_temp_shift_data_reg_41_ ( .D(R2_n172), .CK(clk), .Q(
        R2_U16_DATA1_41) );
  DLH_X1 R2_mix_in_data_reg_40_ ( .G(R2_n2392), .D(R2_U16_DATA1_40), .Q(
        R2_n1169) );
  DFF_X1 R2_temp_shift_data_reg_40_ ( .D(R2_n171), .CK(clk), .Q(
        R2_U16_DATA1_40) );
  DLH_X1 R2_mix_in_data_reg_39_ ( .G(R2_n2393), .D(R2_U16_DATA1_39), .Q(
        R2_n1168) );
  DFF_X1 R2_temp_shift_data_reg_39_ ( .D(R2_n170), .CK(clk), .Q(
        R2_U16_DATA1_39) );
  DLH_X1 R2_mix_in_data_reg_38_ ( .G(R2_n2393), .D(R2_U16_DATA1_38), .Q(
        R2_n1167) );
  DFF_X1 R2_temp_shift_data_reg_38_ ( .D(R2_n169), .CK(clk), .Q(
        R2_U16_DATA1_38) );
  DLH_X1 R2_mix_in_data_reg_37_ ( .G(R2_n2393), .D(R2_U16_DATA1_37), .Q(
        R2_n1166) );
  DFF_X1 R2_temp_shift_data_reg_37_ ( .D(R2_n168), .CK(clk), .Q(
        R2_U16_DATA1_37) );
  DLH_X1 R2_mix_in_data_reg_36_ ( .G(R2_n2393), .D(R2_U16_DATA1_36), .Q(
        R2_n1165) );
  DFF_X1 R2_temp_shift_data_reg_36_ ( .D(R2_n167), .CK(clk), .Q(
        R2_U16_DATA1_36) );
  DLH_X1 R2_mix_in_data_reg_35_ ( .G(R2_n2393), .D(R2_U16_DATA1_35), .Q(
        R2_n1164) );
  DFF_X1 R2_temp_shift_data_reg_35_ ( .D(R2_n166), .CK(clk), .Q(
        R2_U16_DATA1_35) );
  DLH_X1 R2_mix_in_data_reg_34_ ( .G(R2_n2393), .D(R2_U16_DATA1_34), .Q(
        R2_n1163) );
  DFF_X1 R2_temp_shift_data_reg_34_ ( .D(R2_n165), .CK(clk), .Q(
        R2_U16_DATA1_34) );
  DLH_X1 R2_mix_in_data_reg_33_ ( .G(R2_n2393), .D(R2_U16_DATA1_33), .Q(
        R2_n1162) );
  DFF_X1 R2_temp_shift_data_reg_33_ ( .D(R2_n164), .CK(clk), .Q(
        R2_U16_DATA1_33) );
  DLH_X1 R2_mix_in_data_reg_32_ ( .G(R2_n2393), .D(R2_U16_DATA1_32), .Q(
        R2_n1161) );
  DFF_X1 R2_temp_shift_data_reg_32_ ( .D(R2_n163), .CK(clk), .Q(
        R2_U16_DATA1_32) );
  DLH_X1 R2_mix_in_data_reg_31_ ( .G(R2_n2393), .D(R2_U16_DATA1_31), .Q(
        R2_n1160) );
  DFF_X1 R2_temp_shift_data_reg_31_ ( .D(R2_n162), .CK(clk), .Q(
        R2_U16_DATA1_31) );
  DLH_X1 R2_mix_in_data_reg_30_ ( .G(R2_n2393), .D(R2_U16_DATA1_30), .Q(
        R2_n1159) );
  DFF_X1 R2_temp_shift_data_reg_30_ ( .D(R2_n161), .CK(clk), .Q(
        R2_U16_DATA1_30) );
  DLH_X1 R2_mix_in_data_reg_29_ ( .G(R2_n2393), .D(R2_U16_DATA1_29), .Q(
        R2_n1158) );
  DFF_X1 R2_temp_shift_data_reg_29_ ( .D(R2_n160), .CK(clk), .Q(
        R2_U16_DATA1_29) );
  DLH_X1 R2_mix_in_data_reg_28_ ( .G(R2_n2394), .D(R2_U16_DATA1_28), .Q(
        R2_n1157) );
  DFF_X1 R2_temp_shift_data_reg_28_ ( .D(R2_n159), .CK(clk), .Q(
        R2_U16_DATA1_28) );
  DLH_X1 R2_mix_in_data_reg_27_ ( .G(R2_n2392), .D(R2_U16_DATA1_27), .Q(
        R2_n1156) );
  DFF_X1 R2_temp_shift_data_reg_27_ ( .D(R2_n158), .CK(clk), .Q(
        R2_U16_DATA1_27) );
  DLH_X1 R2_mix_in_data_reg_26_ ( .G(R2_n2394), .D(R2_U16_DATA1_26), .Q(
        R2_n1155) );
  DFF_X1 R2_temp_shift_data_reg_26_ ( .D(R2_n157), .CK(clk), .Q(
        R2_U16_DATA1_26) );
  DLH_X1 R2_mix_in_data_reg_25_ ( .G(R2_n2392), .D(R2_U16_DATA1_25), .Q(
        R2_n1154) );
  DFF_X1 R2_temp_shift_data_reg_25_ ( .D(R2_n156), .CK(clk), .Q(
        R2_U16_DATA1_25) );
  DLH_X1 R2_mix_in_data_reg_24_ ( .G(R2_n2391), .D(R2_U16_DATA1_24), .Q(
        R2_n1153) );
  DFF_X1 R2_temp_shift_data_reg_24_ ( .D(R2_n155), .CK(clk), .Q(
        R2_U16_DATA1_24) );
  DLH_X1 R2_mix_in_data_reg_23_ ( .G(R2_n2391), .D(R2_U16_DATA1_23), .Q(
        R2_n1152) );
  DFF_X1 R2_temp_shift_data_reg_23_ ( .D(R2_n154), .CK(clk), .Q(
        R2_U16_DATA1_23) );
  DLH_X1 R2_mix_in_data_reg_22_ ( .G(R2_n2394), .D(R2_U16_DATA1_22), .Q(
        R2_n1151) );
  DFF_X1 R2_temp_shift_data_reg_22_ ( .D(R2_n153), .CK(clk), .Q(
        R2_U16_DATA1_22) );
  DLH_X1 R2_mix_in_data_reg_21_ ( .G(R2_n2394), .D(R2_U16_DATA1_21), .Q(
        R2_n1150) );
  DFF_X1 R2_temp_shift_data_reg_21_ ( .D(R2_n152), .CK(clk), .Q(
        R2_U16_DATA1_21) );
  DLH_X1 R2_mix_in_data_reg_20_ ( .G(R2_n2392), .D(R2_U16_DATA1_20), .Q(
        R2_n1149) );
  DFF_X1 R2_temp_shift_data_reg_20_ ( .D(R2_n151), .CK(clk), .Q(
        R2_U16_DATA1_20) );
  DLH_X1 R2_mix_in_data_reg_19_ ( .G(R2_n2392), .D(R2_U16_DATA1_19), .Q(
        R2_n1148) );
  DFF_X1 R2_temp_shift_data_reg_19_ ( .D(R2_n150), .CK(clk), .Q(
        R2_U16_DATA1_19) );
  DLH_X1 R2_mix_in_data_reg_18_ ( .G(R2_n2392), .D(R2_U16_DATA1_18), .Q(
        R2_n1147) );
  DFF_X1 R2_temp_shift_data_reg_18_ ( .D(R2_n149), .CK(clk), .Q(
        R2_U16_DATA1_18) );
  DLH_X1 R2_mix_in_data_reg_17_ ( .G(R2_n2394), .D(R2_U16_DATA1_17), .Q(
        R2_n1146) );
  DFF_X1 R2_temp_shift_data_reg_17_ ( .D(R2_n148), .CK(clk), .Q(
        R2_U16_DATA1_17) );
  DLH_X1 R2_mix_in_data_reg_16_ ( .G(R2_n2394), .D(R2_U16_DATA1_16), .Q(
        R2_n1145) );
  DFF_X1 R2_temp_shift_data_reg_16_ ( .D(R2_n147), .CK(clk), .Q(
        R2_U16_DATA1_16) );
  DLH_X1 R2_mix_in_data_reg_15_ ( .G(R2_n2394), .D(R2_U16_DATA1_15), .Q(
        R2_n1144) );
  DFF_X1 R2_temp_shift_data_reg_15_ ( .D(R2_n146), .CK(clk), .Q(
        R2_U16_DATA1_15) );
  DLH_X1 R2_mix_in_data_reg_14_ ( .G(R2_n2394), .D(R2_U16_DATA1_14), .Q(
        R2_n1143) );
  DFF_X1 R2_temp_shift_data_reg_14_ ( .D(R2_n145), .CK(clk), .Q(
        R2_U16_DATA1_14) );
  DLH_X1 R2_mix_in_data_reg_13_ ( .G(R2_n2394), .D(R2_U16_DATA1_13), .Q(
        R2_n1142) );
  DFF_X1 R2_temp_shift_data_reg_13_ ( .D(R2_n144), .CK(clk), .Q(
        R2_U16_DATA1_13) );
  DLH_X1 R2_mix_in_data_reg_12_ ( .G(R2_n2394), .D(R2_U16_DATA1_12), .Q(
        R2_n1141) );
  DFF_X1 R2_temp_shift_data_reg_12_ ( .D(R2_n143), .CK(clk), .Q(
        R2_U16_DATA1_12) );
  DLH_X1 R2_mix_in_data_reg_11_ ( .G(R2_n2394), .D(R2_U16_DATA1_11), .Q(
        R2_n1140) );
  DFF_X1 R2_temp_shift_data_reg_11_ ( .D(R2_n142), .CK(clk), .Q(
        R2_U16_DATA1_11) );
  DLH_X1 R2_mix_in_data_reg_10_ ( .G(R2_n2394), .D(R2_U16_DATA1_10), .Q(
        R2_n1139) );
  DFF_X1 R2_temp_shift_data_reg_10_ ( .D(R2_n141), .CK(clk), .Q(
        R2_U16_DATA1_10) );
  DLH_X1 R2_mix_in_data_reg_9_ ( .G(R2_n2394), .D(R2_U16_DATA1_9), .Q(R2_n1138) );
  DFF_X1 R2_temp_shift_data_reg_9_ ( .D(R2_n140), .CK(clk), .Q(R2_U16_DATA1_9)
         );
  DLH_X1 R2_mix_in_data_reg_8_ ( .G(R2_n2394), .D(R2_U16_DATA1_8), .Q(R2_n1137) );
  DFF_X1 R2_temp_shift_data_reg_8_ ( .D(R2_n139), .CK(clk), .Q(R2_U16_DATA1_8)
         );
  DLH_X1 R2_mix_in_data_reg_7_ ( .G(R2_n2394), .D(R2_U16_DATA1_7), .Q(R2_n1136) );
  DFF_X1 R2_temp_shift_data_reg_7_ ( .D(R2_n138), .CK(clk), .Q(R2_U16_DATA1_7)
         );
  DLH_X1 R2_mix_in_data_reg_6_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_6), .Q(
        R2_n1135) );
  DFF_X1 R2_temp_shift_data_reg_6_ ( .D(R2_n137), .CK(clk), .Q(R2_U16_DATA1_6)
         );
  DLH_X1 R2_mix_in_data_reg_5_ ( .G(R2_n2393), .D(R2_U16_DATA1_5), .Q(R2_n1134) );
  DFF_X1 R2_temp_shift_data_reg_5_ ( .D(R2_n136), .CK(clk), .Q(R2_U16_DATA1_5)
         );
  DLH_X1 R2_mix_in_data_reg_4_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_4), .Q(
        R2_n1133) );
  DFF_X1 R2_temp_shift_data_reg_4_ ( .D(R2_n135), .CK(clk), .Q(R2_U16_DATA1_4)
         );
  DLH_X1 R2_mix_in_data_reg_3_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_3), .Q(
        R2_n1132) );
  DFF_X1 R2_temp_shift_data_reg_3_ ( .D(R2_n134), .CK(clk), .Q(R2_U16_DATA1_3)
         );
  DLH_X1 R2_mix_in_data_reg_2_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_2), .Q(
        R2_n1131) );
  DFF_X1 R2_temp_shift_data_reg_2_ ( .D(R2_n133), .CK(clk), .Q(R2_U16_DATA1_2)
         );
  DLH_X1 R2_mix_in_data_reg_1_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_1), .Q(
        R2_n1130) );
  DFF_X1 R2_temp_shift_data_reg_1_ ( .D(R2_n132), .CK(clk), .Q(R2_U16_DATA1_1)
         );
  DLH_X1 R2_mix_in_data_reg_0_ ( .G(R2_U21_Z_1), .D(R2_U16_DATA1_0), .Q(
        R2_n1129) );
  DFF_X1 R2_temp_shift_data_reg_0_ ( .D(R2_n131), .CK(clk), .Q(R2_U16_DATA1_0)
         );
  DLH_X1 R2_add_key_in_reg_70_ ( .G(R2_n2402), .D(n3462), .Q(R2_n814) );
  DLH_X1 R2_add_key_in_reg_71_ ( .G(R2_U23_Z_1), .D(n3463), .Q(R2_n815) );
  DLH_X1 R2_add_key_in_reg_72_ ( .G(R2_n2400), .D(n3464), .Q(R2_n816) );
  DLH_X1 R2_add_key_in_reg_73_ ( .G(R2_n2403), .D(n3465), .Q(R2_n817) );
  DLH_X1 R2_add_key_in_reg_74_ ( .G(R2_n2400), .D(n3466), .Q(R2_n818) );
  DLH_X1 R2_add_key_in_reg_75_ ( .G(R2_n2401), .D(n3467), .Q(R2_n819) );
  DLH_X1 R2_add_key_in_reg_76_ ( .G(R2_n2401), .D(n3468), .Q(R2_n820) );
  DLH_X1 R2_add_key_in_reg_77_ ( .G(R2_n2404), .D(n3469), .Q(R2_n821) );
  DLH_X1 R2_add_key_in_reg_78_ ( .G(R2_n2404), .D(n3470), .Q(R2_n822) );
  DLH_X1 R2_add_key_in_reg_79_ ( .G(R2_n2400), .D(n3471), .Q(R2_n823) );
  DLH_X1 R2_add_key_in_reg_80_ ( .G(R2_U23_Z_1), .D(n3472), .Q(R2_n824) );
  DLH_X1 R2_add_key_in_reg_81_ ( .G(R2_n2401), .D(n3473), .Q(R2_n825) );
  DLH_X1 R2_add_key_in_reg_82_ ( .G(R2_n2398), .D(n3474), .Q(R2_n826) );
  DLH_X1 R2_add_key_in_reg_83_ ( .G(R2_n2401), .D(n3475), .Q(R2_n827) );
  DLH_X1 R2_add_key_in_reg_84_ ( .G(R2_n2403), .D(n3476), .Q(R2_n828) );
  DLH_X1 R2_add_key_in_reg_85_ ( .G(R2_n2399), .D(n3477), .Q(R2_n829) );
  DLH_X1 R2_add_key_in_reg_86_ ( .G(R2_n2398), .D(n3478), .Q(R2_n830) );
  DLH_X1 R2_add_key_in_reg_87_ ( .G(R2_n2398), .D(n3479), .Q(R2_n831) );
  DLH_X1 R2_add_key_in_reg_88_ ( .G(R2_n2401), .D(n3480), .Q(R2_n832) );
  DLH_X1 R2_add_key_in_reg_89_ ( .G(R2_U23_Z_1), .D(n3481), .Q(R2_n833) );
  DLH_X1 R2_add_key_in_reg_90_ ( .G(R2_n2404), .D(n3482), .Q(R2_n834) );
  DLH_X1 R2_add_key_in_reg_91_ ( .G(R2_n2398), .D(n3483), .Q(R2_n835) );
  DLH_X1 R2_add_key_in_reg_92_ ( .G(R2_n2400), .D(n3484), .Q(R2_n836) );
  DLH_X1 R2_add_key_in_reg_93_ ( .G(R2_U23_Z_1), .D(n3485), .Q(R2_n837) );
  DLH_X1 R2_add_key_in_reg_94_ ( .G(R2_n2402), .D(n3486), .Q(R2_n838) );
  DLH_X1 R2_add_key_in_reg_95_ ( .G(R2_n2401), .D(n3487), .Q(R2_n839) );
  DLH_X1 R2_add_key_in_reg_96_ ( .G(R2_n2399), .D(n3488), .Q(R2_n840) );
  DLH_X1 R2_add_key_in_reg_97_ ( .G(R2_n2399), .D(n3489), .Q(R2_n841) );
  DLH_X1 R2_add_key_in_reg_98_ ( .G(R2_n2399), .D(n3490), .Q(R2_n842) );
  DLH_X1 R2_add_key_in_reg_99_ ( .G(R2_n2399), .D(n3491), .Q(R2_n843) );
  DLH_X1 R2_add_key_in_reg_100_ ( .G(R2_n2399), .D(n3492), .Q(R2_n844) );
  DLH_X1 R2_add_key_in_reg_101_ ( .G(R2_n2399), .D(n3493), .Q(R2_n845) );
  DLH_X1 R2_add_key_in_reg_102_ ( .G(R2_n2399), .D(n3494), .Q(R2_n846) );
  DLH_X1 R2_add_key_in_reg_103_ ( .G(R2_n2399), .D(n3495), .Q(R2_n847) );
  DLH_X1 R2_add_key_in_reg_104_ ( .G(R2_n2399), .D(n3496), .Q(R2_n848) );
  DLH_X1 R2_add_key_in_reg_105_ ( .G(R2_n2399), .D(n3497), .Q(R2_n849) );
  DLH_X1 R2_add_key_in_reg_106_ ( .G(R2_n2399), .D(n3498), .Q(R2_n850) );
  DLH_X1 R2_add_key_in_reg_107_ ( .G(R2_n2400), .D(n3499), .Q(R2_n851) );
  DLH_X1 R2_add_key_in_reg_108_ ( .G(R2_n2402), .D(n3500), .Q(R2_n852) );
  DLH_X1 R2_add_key_in_reg_109_ ( .G(R2_n2404), .D(n3501), .Q(R2_n853) );
  DLH_X1 R2_add_key_in_reg_110_ ( .G(R2_n2403), .D(n3502), .Q(R2_n854) );
  DLH_X1 R2_add_key_in_reg_111_ ( .G(R2_n2404), .D(n3503), .Q(R2_n855) );
  DLH_X1 R2_add_key_in_reg_112_ ( .G(R2_n2404), .D(n3504), .Q(R2_n856) );
  DLH_X1 R2_add_key_in_reg_113_ ( .G(R2_n2398), .D(n3505), .Q(R2_n857) );
  DLH_X1 R2_add_key_in_reg_114_ ( .G(R2_n2403), .D(n3506), .Q(R2_n858) );
  DLH_X1 R2_add_key_in_reg_115_ ( .G(R2_n2399), .D(n3507), .Q(R2_n859) );
  DLH_X1 R2_add_key_in_reg_116_ ( .G(R2_n2403), .D(n3508), .Q(R2_n860) );
  DLH_X1 R2_add_key_in_reg_117_ ( .G(R2_U23_Z_1), .D(n3509), .Q(R2_n861) );
  DLH_X1 R2_add_key_in_reg_118_ ( .G(R2_n2398), .D(n3510), .Q(R2_n862) );
  DLH_X1 R2_add_key_in_reg_119_ ( .G(R2_n2403), .D(n3511), .Q(R2_n863) );
  DLH_X1 R2_add_key_in_reg_120_ ( .G(R2_n2399), .D(n3512), .Q(R2_n864) );
  DLH_X1 R2_add_key_in_reg_121_ ( .G(R2_n2401), .D(n3513), .Q(R2_n865) );
  DLH_X1 R2_add_key_in_reg_122_ ( .G(R2_n2403), .D(n3514), .Q(R2_n866) );
  DLH_X1 R2_add_key_in_reg_123_ ( .G(R2_n2400), .D(n3515), .Q(R2_n867) );
  DLH_X1 R2_add_key_in_reg_124_ ( .G(R2_U23_Z_1), .D(n3516), .Q(R2_n868) );
  DLH_X1 R2_add_key_in_reg_125_ ( .G(R2_n2399), .D(n3517), .Q(R2_n869) );
  DLH_X1 R2_add_key_in_reg_126_ ( .G(R2_n2404), .D(n3518), .Q(R2_n870) );
  DLH_X1 R2_add_key_in_reg_127_ ( .G(R2_n2402), .D(n3519), .Q(R2_n871) );
  DLH_X1 R2_add_key_in_reg_0_ ( .G(R2_n2399), .D(n3392), .Q(R2_n744) );
  DLH_X1 R2_add_key_in_reg_1_ ( .G(R2_n2400), .D(n3393), .Q(R2_n745) );
  DLH_X1 R2_add_key_in_reg_2_ ( .G(R2_n2400), .D(n3394), .Q(R2_n746) );
  DLH_X1 R2_add_key_in_reg_3_ ( .G(R2_n2400), .D(n3395), .Q(R2_n747) );
  DLH_X1 R2_add_key_in_reg_4_ ( .G(R2_n2400), .D(n3396), .Q(R2_n748) );
  DLH_X1 R2_add_key_in_reg_5_ ( .G(R2_n2400), .D(n3397), .Q(R2_n749) );
  DLH_X1 R2_add_key_in_reg_6_ ( .G(R2_n2400), .D(n3398), .Q(R2_n750) );
  DLH_X1 R2_add_key_in_reg_7_ ( .G(R2_n2400), .D(n3399), .Q(R2_n751) );
  DLH_X1 R2_add_key_in_reg_8_ ( .G(R2_n2400), .D(n3400), .Q(R2_n752) );
  DLH_X1 R2_add_key_in_reg_9_ ( .G(R2_n2400), .D(n3401), .Q(R2_n753) );
  DLH_X1 R2_add_key_in_reg_10_ ( .G(R2_n2400), .D(n3402), .Q(R2_n754) );
  DLH_X1 R2_add_key_in_reg_11_ ( .G(R2_n2400), .D(n3403), .Q(R2_n755) );
  DLH_X1 R2_add_key_in_reg_12_ ( .G(R2_n2398), .D(n3404), .Q(R2_n756) );
  DLH_X1 R2_add_key_in_reg_13_ ( .G(R2_n2400), .D(n3405), .Q(R2_n757) );
  DLH_X1 R2_add_key_in_reg_14_ ( .G(R2_n2400), .D(n3406), .Q(R2_n758) );
  DLH_X1 R2_add_key_in_reg_15_ ( .G(R2_n2404), .D(n3407), .Q(R2_n759) );
  DLH_X1 R2_add_key_in_reg_16_ ( .G(R2_n2401), .D(n3408), .Q(R2_n760) );
  DLH_X1 R2_add_key_in_reg_17_ ( .G(R2_n2402), .D(n3409), .Q(R2_n761) );
  DLH_X1 R2_add_key_in_reg_18_ ( .G(R2_n2404), .D(n3410), .Q(R2_n762) );
  DLH_X1 R2_add_key_in_reg_19_ ( .G(R2_n2403), .D(n3411), .Q(R2_n763) );
  DLH_X1 R2_add_key_in_reg_20_ ( .G(R2_n2402), .D(n3412), .Q(R2_n764) );
  DLH_X1 R2_add_key_in_reg_21_ ( .G(R2_n2402), .D(n3413), .Q(R2_n765) );
  DLH_X1 R2_add_key_in_reg_22_ ( .G(R2_n2399), .D(n3414), .Q(R2_n766) );
  DLH_X1 R2_add_key_in_reg_23_ ( .G(R2_n2402), .D(n3415), .Q(R2_n767) );
  DLH_X1 R2_add_key_in_reg_24_ ( .G(R2_n2402), .D(n3416), .Q(R2_n768) );
  DLH_X1 R2_add_key_in_reg_25_ ( .G(R2_n2403), .D(n3417), .Q(R2_n769) );
  DLH_X1 R2_add_key_in_reg_26_ ( .G(R2_n2403), .D(n3418), .Q(R2_n770) );
  DLH_X1 R2_add_key_in_reg_27_ ( .G(R2_n2404), .D(n3419), .Q(R2_n771) );
  DLH_X1 R2_add_key_in_reg_28_ ( .G(R2_n2403), .D(n3420), .Q(R2_n772) );
  DLH_X1 R2_add_key_in_reg_29_ ( .G(R2_n2401), .D(n3421), .Q(R2_n773) );
  DLH_X1 R2_add_key_in_reg_30_ ( .G(R2_n2401), .D(n3422), .Q(R2_n774) );
  DLH_X1 R2_add_key_in_reg_31_ ( .G(R2_n2403), .D(n3423), .Q(R2_n775) );
  DLH_X1 R2_add_key_in_reg_32_ ( .G(R2_n2404), .D(n3424), .Q(R2_n776) );
  DLH_X1 R2_add_key_in_reg_33_ ( .G(R2_n2402), .D(n3425), .Q(R2_n777) );
  DLH_X1 R2_add_key_in_reg_34_ ( .G(R2_n2402), .D(n3426), .Q(R2_n778) );
  DLH_X1 R2_add_key_in_reg_35_ ( .G(R2_n2404), .D(n3427), .Q(R2_n779) );
  DLH_X1 R2_add_key_in_reg_36_ ( .G(R2_n2404), .D(n3428), .Q(R2_n780) );
  DLH_X1 R2_add_key_in_reg_37_ ( .G(R2_n2401), .D(n3429), .Q(R2_n781) );
  DLH_X1 R2_add_key_in_reg_38_ ( .G(R2_n2401), .D(n3430), .Q(R2_n782) );
  DLH_X1 R2_add_key_in_reg_39_ ( .G(R2_n2403), .D(n3431), .Q(R2_n783) );
  DLH_X1 R2_add_key_in_reg_40_ ( .G(R2_n2401), .D(n3432), .Q(R2_n784) );
  DLH_X1 R2_add_key_in_reg_41_ ( .G(R2_n2404), .D(n3433), .Q(R2_n785) );
  DLH_X1 R2_add_key_in_reg_42_ ( .G(R2_n2403), .D(n3434), .Q(R2_n786) );
  DLH_X1 R2_add_key_in_reg_43_ ( .G(R2_n2402), .D(n3435), .Q(R2_n787) );
  DLH_X1 R2_add_key_in_reg_44_ ( .G(R2_n2401), .D(n3436), .Q(R2_n788) );
  DLH_X1 R2_add_key_in_reg_45_ ( .G(R2_n2402), .D(n3437), .Q(R2_n789) );
  DLH_X1 R2_add_key_in_reg_46_ ( .G(R2_n2401), .D(n3438), .Q(R2_n790) );
  DLH_X1 R2_add_key_in_reg_47_ ( .G(R2_n2403), .D(n3439), .Q(R2_n791) );
  DLH_X1 R2_add_key_in_reg_48_ ( .G(R2_n2398), .D(n3440), .Q(R2_n792) );
  DLH_X1 R2_add_key_in_reg_49_ ( .G(R2_U23_Z_1), .D(n3441), .Q(R2_n793) );
  DLH_X1 R2_add_key_in_reg_50_ ( .G(R2_U23_Z_1), .D(n3442), .Q(R2_n794) );
  DLH_X1 R2_add_key_in_reg_51_ ( .G(R2_n2402), .D(n3443), .Q(R2_n795) );
  DLH_X1 R2_add_key_in_reg_52_ ( .G(R2_n2400), .D(n3444), .Q(R2_n796) );
  DLH_X1 R2_add_key_in_reg_53_ ( .G(R2_n2399), .D(n3445), .Q(R2_n797) );
  DLH_X1 R2_add_key_in_reg_54_ ( .G(R2_n2403), .D(n3446), .Q(R2_n798) );
  DLH_X1 R2_add_key_in_reg_55_ ( .G(R2_n2404), .D(n3447), .Q(R2_n799) );
  DLH_X1 R2_add_key_in_reg_56_ ( .G(R2_n2401), .D(n3448), .Q(R2_n800) );
  DLH_X1 R2_add_key_in_reg_57_ ( .G(R2_n2402), .D(n3449), .Q(R2_n801) );
  DLH_X1 R2_add_key_in_reg_58_ ( .G(R2_n2403), .D(n3450), .Q(R2_n802) );
  DLH_X1 R2_add_key_in_reg_59_ ( .G(R2_n2404), .D(n3451), .Q(R2_n803) );
  DLH_X1 R2_add_key_in_reg_60_ ( .G(R2_n2401), .D(n3452), .Q(R2_n804) );
  DLH_X1 R2_add_key_in_reg_61_ ( .G(R2_n2403), .D(n3453), .Q(R2_n805) );
  DLH_X1 R2_add_key_in_reg_62_ ( .G(R2_n2402), .D(n3454), .Q(R2_n806) );
  DLH_X1 R2_add_key_in_reg_63_ ( .G(R2_n2402), .D(n3455), .Q(R2_n807) );
  DLH_X1 R2_add_key_in_reg_64_ ( .G(R2_n2403), .D(n3456), .Q(R2_n808) );
  DLH_X1 R2_add_key_in_reg_65_ ( .G(R2_n2404), .D(n3457), .Q(R2_n809) );
  DLH_X1 R2_add_key_in_reg_66_ ( .G(R2_n2402), .D(n3458), .Q(R2_n810) );
  DLH_X1 R2_add_key_in_reg_67_ ( .G(R2_n2404), .D(n3459), .Q(R2_n811) );
  DLH_X1 R2_add_key_in_reg_68_ ( .G(R2_n2401), .D(n3460), .Q(R2_n812) );
  DLH_X1 R2_add_key_in_reg_69_ ( .G(R2_n2402), .D(n3461), .Q(R2_n813) );
  DLH_X1 R2_shift_in_data_reg_98_ ( .G(R2_n2397), .D(R2_n580), .Q(R2_n1484) );
  DLH_X1 R2_shift_in_data_reg_97_ ( .G(R2_U22_Z_1), .D(R2_n579), .Q(R2_n1483)
         );
  DLH_X1 R2_shift_in_data_reg_96_ ( .G(R2_U22_Z_1), .D(R2_n578), .Q(R2_n1482)
         );
  DLH_X1 R2_shift_in_data_reg_95_ ( .G(R2_U22_Z_1), .D(R2_n577), .Q(R2_n1481)
         );
  DLH_X1 R2_shift_in_data_reg_94_ ( .G(R2_n2395), .D(R2_n576), .Q(R2_n1480) );
  DLH_X1 R2_shift_in_data_reg_93_ ( .G(R2_U22_Z_1), .D(R2_n575), .Q(R2_n1479)
         );
  DLH_X1 R2_shift_in_data_reg_92_ ( .G(R2_n2395), .D(R2_n574), .Q(R2_n1478) );
  DLH_X1 R2_shift_in_data_reg_91_ ( .G(R2_n2395), .D(R2_n573), .Q(R2_n1477) );
  DLH_X1 R2_shift_in_data_reg_90_ ( .G(R2_U22_Z_1), .D(R2_n572), .Q(R2_n1476)
         );
  DLH_X1 R2_shift_in_data_reg_89_ ( .G(R2_U22_Z_1), .D(R2_n571), .Q(R2_n1475)
         );
  DLH_X1 R2_shift_in_data_reg_88_ ( .G(R2_n2397), .D(R2_n570), .Q(R2_n1474) );
  DLH_X1 R2_shift_in_data_reg_87_ ( .G(R2_n2397), .D(R2_n569), .Q(R2_n1473) );
  DLH_X1 R2_shift_in_data_reg_86_ ( .G(R2_U22_Z_1), .D(R2_n568), .Q(R2_n1472)
         );
  DLH_X1 R2_shift_in_data_reg_85_ ( .G(R2_n2397), .D(R2_n567), .Q(R2_n1471) );
  DLH_X1 R2_shift_in_data_reg_84_ ( .G(R2_n2396), .D(R2_n566), .Q(R2_n1470) );
  DLH_X1 R2_shift_in_data_reg_83_ ( .G(R2_n2395), .D(R2_n565), .Q(R2_n1469) );
  DLH_X1 R2_shift_in_data_reg_82_ ( .G(R2_U22_Z_1), .D(R2_n564), .Q(R2_n1468)
         );
  DLH_X1 R2_shift_in_data_reg_81_ ( .G(R2_n2396), .D(R2_n563), .Q(R2_n1467) );
  DLH_X1 R2_shift_in_data_reg_80_ ( .G(R2_U22_Z_1), .D(R2_n562), .Q(R2_n1466)
         );
  DLH_X1 R2_shift_in_data_reg_79_ ( .G(R2_n2397), .D(R2_n561), .Q(R2_n1465) );
  DLH_X1 R2_shift_in_data_reg_78_ ( .G(R2_n2395), .D(R2_n560), .Q(R2_n1464) );
  DLH_X1 R2_shift_in_data_reg_77_ ( .G(R2_n2395), .D(R2_n559), .Q(R2_n1463) );
  DLH_X1 R2_shift_in_data_reg_76_ ( .G(R2_n2397), .D(R2_n558), .Q(R2_n1462) );
  DLH_X1 R2_shift_in_data_reg_75_ ( .G(R2_n2396), .D(R2_n557), .Q(R2_n1461) );
  DLH_X1 R2_shift_in_data_reg_74_ ( .G(R2_U22_Z_1), .D(R2_n556), .Q(R2_n1460)
         );
  DLH_X1 R2_shift_in_data_reg_73_ ( .G(R2_n2395), .D(R2_n555), .Q(R2_n1459) );
  DLH_X1 R2_shift_in_data_reg_72_ ( .G(R2_n2396), .D(R2_n554), .Q(R2_n1458) );
  DLH_X1 R2_shift_in_data_reg_71_ ( .G(R2_U22_Z_1), .D(R2_n553), .Q(R2_n1457)
         );
  DLH_X1 R2_shift_in_data_reg_70_ ( .G(R2_n2397), .D(R2_n552), .Q(R2_n1456) );
  DLH_X1 R2_shift_in_data_reg_69_ ( .G(R2_n2395), .D(R2_n551), .Q(R2_n1455) );
  DLH_X1 R2_shift_in_data_reg_68_ ( .G(R2_U22_Z_1), .D(R2_n550), .Q(R2_n1454)
         );
  DLH_X1 R2_shift_in_data_reg_67_ ( .G(R2_U22_Z_1), .D(R2_n549), .Q(R2_n1453)
         );
  DLH_X1 R2_shift_in_data_reg_66_ ( .G(R2_n2395), .D(R2_n548), .Q(R2_n1452) );
  DLH_X1 R2_shift_in_data_reg_65_ ( .G(R2_n2397), .D(R2_n547), .Q(R2_n1451) );
  DLH_X1 R2_shift_in_data_reg_64_ ( .G(R2_n2396), .D(R2_n546), .Q(R2_n1450) );
  DLH_X1 R2_shift_in_data_reg_63_ ( .G(R2_n2397), .D(R2_n545), .Q(R2_n1449) );
  DLH_X1 R2_shift_in_data_reg_62_ ( .G(R2_n2396), .D(R2_n544), .Q(R2_n1448) );
  DLH_X1 R2_shift_in_data_reg_61_ ( .G(R2_n2395), .D(R2_n543), .Q(R2_n1447) );
  DLH_X1 R2_shift_in_data_reg_60_ ( .G(R2_n2395), .D(R2_n542), .Q(R2_n1446) );
  DLH_X1 R2_shift_in_data_reg_59_ ( .G(R2_U22_Z_1), .D(R2_n541), .Q(R2_n1445)
         );
  DLH_X1 R2_shift_in_data_reg_58_ ( .G(R2_n2397), .D(R2_n540), .Q(R2_n1444) );
  DLH_X1 R2_shift_in_data_reg_57_ ( .G(R2_n2396), .D(R2_n539), .Q(R2_n1443) );
  DLH_X1 R2_shift_in_data_reg_56_ ( .G(R2_n2396), .D(R2_n538), .Q(R2_n1442) );
  DLH_X1 R2_shift_in_data_reg_55_ ( .G(R2_n2396), .D(R2_n537), .Q(R2_n1441) );
  DLH_X1 R2_shift_in_data_reg_54_ ( .G(R2_n2395), .D(R2_n536), .Q(R2_n1440) );
  DLH_X1 R2_shift_in_data_reg_53_ ( .G(R2_U22_Z_1), .D(R2_n535), .Q(R2_n1439)
         );
  DLH_X1 R2_shift_in_data_reg_52_ ( .G(R2_n2397), .D(R2_n534), .Q(R2_n1438) );
  DLH_X1 R2_shift_in_data_reg_51_ ( .G(R2_U22_Z_1), .D(R2_n533), .Q(R2_n1437)
         );
  DLH_X1 R2_shift_in_data_reg_50_ ( .G(R2_U22_Z_1), .D(R2_n532), .Q(R2_n1436)
         );
  DLH_X1 R2_shift_in_data_reg_49_ ( .G(R2_n2396), .D(R2_n531), .Q(R2_n1435) );
  DLH_X1 R2_shift_in_data_reg_48_ ( .G(R2_n2397), .D(R2_n530), .Q(R2_n1434) );
  DLH_X1 R2_shift_in_data_reg_47_ ( .G(R2_n2397), .D(R2_n529), .Q(R2_n1433) );
  DLH_X1 R2_shift_in_data_reg_46_ ( .G(R2_n2397), .D(R2_n528), .Q(R2_n1432) );
  DLH_X1 R2_shift_in_data_reg_45_ ( .G(R2_n2395), .D(R2_n527), .Q(R2_n1431) );
  DLH_X1 R2_shift_in_data_reg_44_ ( .G(R2_n2396), .D(R2_n526), .Q(R2_n1430) );
  DLH_X1 R2_shift_in_data_reg_43_ ( .G(R2_n2395), .D(R2_n525), .Q(R2_n1429) );
  DLH_X1 R2_shift_in_data_reg_42_ ( .G(R2_U22_Z_1), .D(R2_n524), .Q(R2_n1428)
         );
  DLH_X1 R2_shift_in_data_reg_41_ ( .G(R2_U22_Z_1), .D(R2_n523), .Q(R2_n1427)
         );
  DLH_X1 R2_shift_in_data_reg_40_ ( .G(R2_n2395), .D(R2_n522), .Q(R2_n1426) );
  DLH_X1 R2_shift_in_data_reg_39_ ( .G(R2_n2396), .D(R2_n521), .Q(R2_n1425) );
  DLH_X1 R2_shift_in_data_reg_38_ ( .G(R2_U22_Z_1), .D(R2_n520), .Q(R2_n1424)
         );
  DLH_X1 R2_shift_in_data_reg_37_ ( .G(R2_n2397), .D(R2_n519), .Q(R2_n1423) );
  DLH_X1 R2_shift_in_data_reg_36_ ( .G(R2_n2395), .D(R2_n518), .Q(R2_n1422) );
  DLH_X1 R2_shift_in_data_reg_35_ ( .G(R2_n2395), .D(R2_n517), .Q(R2_n1421) );
  DLH_X1 R2_shift_in_data_reg_34_ ( .G(R2_U22_Z_1), .D(R2_n516), .Q(R2_n1420)
         );
  DLH_X1 R2_shift_in_data_reg_33_ ( .G(R2_n2395), .D(R2_n515), .Q(R2_n1419) );
  DLH_X1 R2_shift_in_data_reg_32_ ( .G(R2_n2395), .D(R2_n514), .Q(R2_n1418) );
  DLH_X1 R2_shift_in_data_reg_31_ ( .G(R2_n2395), .D(R2_n513), .Q(R2_n1417) );
  DLH_X1 R2_shift_in_data_reg_30_ ( .G(R2_n2396), .D(R2_n512), .Q(R2_n1416) );
  DLH_X1 R2_shift_in_data_reg_29_ ( .G(R2_n2396), .D(R2_n511), .Q(R2_n1415) );
  DLH_X1 R2_shift_in_data_reg_28_ ( .G(R2_n2397), .D(R2_n510), .Q(R2_n1414) );
  DLH_X1 R2_shift_in_data_reg_27_ ( .G(R2_U22_Z_1), .D(R2_n509), .Q(R2_n1413)
         );
  DLH_X1 R2_shift_in_data_reg_26_ ( .G(R2_n2395), .D(R2_n508), .Q(R2_n1412) );
  DLH_X1 R2_shift_in_data_reg_25_ ( .G(R2_n2397), .D(R2_n507), .Q(R2_n1411) );
  DLH_X1 R2_shift_in_data_reg_24_ ( .G(R2_n2395), .D(R2_n506), .Q(R2_n1410) );
  DLH_X1 R2_shift_in_data_reg_23_ ( .G(R2_U22_Z_1), .D(R2_n505), .Q(R2_n1409)
         );
  DLH_X1 R2_shift_in_data_reg_22_ ( .G(R2_n2395), .D(R2_n504), .Q(R2_n1408) );
  DLH_X1 R2_shift_in_data_reg_21_ ( .G(R2_n2397), .D(R2_n503), .Q(R2_n1407) );
  DLH_X1 R2_shift_in_data_reg_20_ ( .G(R2_U22_Z_1), .D(R2_n502), .Q(R2_n1406)
         );
  DLH_X1 R2_shift_in_data_reg_19_ ( .G(R2_n2396), .D(R2_n501), .Q(R2_n1405) );
  DLH_X1 R2_shift_in_data_reg_18_ ( .G(R2_n2395), .D(R2_n500), .Q(R2_n1404) );
  DLH_X1 R2_shift_in_data_reg_17_ ( .G(R2_U22_Z_1), .D(R2_n499), .Q(R2_n1403)
         );
  DLH_X1 R2_shift_in_data_reg_16_ ( .G(R2_n2396), .D(R2_n498), .Q(R2_n1402) );
  DLH_X1 R2_shift_in_data_reg_15_ ( .G(R2_n2396), .D(R2_n497), .Q(R2_n1401) );
  DLH_X1 R2_shift_in_data_reg_14_ ( .G(R2_n2396), .D(R2_n496), .Q(R2_n1400) );
  DLH_X1 R2_shift_in_data_reg_13_ ( .G(R2_n2396), .D(R2_n495), .Q(R2_n1399) );
  DLH_X1 R2_shift_in_data_reg_12_ ( .G(R2_n2397), .D(R2_n494), .Q(R2_n1398) );
  DLH_X1 R2_shift_in_data_reg_11_ ( .G(R2_n2395), .D(R2_n493), .Q(R2_n1397) );
  DLH_X1 R2_shift_in_data_reg_10_ ( .G(R2_U22_Z_1), .D(R2_n492), .Q(R2_n1396)
         );
  DLH_X1 R2_shift_in_data_reg_9_ ( .G(R2_n2396), .D(R2_n491), .Q(R2_n1395) );
  DLH_X1 R2_shift_in_data_reg_8_ ( .G(R2_U22_Z_1), .D(R2_n490), .Q(R2_n1394)
         );
  DLH_X1 R2_shift_in_data_reg_7_ ( .G(R2_n2396), .D(R2_n489), .Q(R2_n1393) );
  DLH_X1 R2_shift_in_data_reg_6_ ( .G(R2_n2396), .D(R2_n488), .Q(R2_n1392) );
  DLH_X1 R2_shift_in_data_reg_5_ ( .G(R2_n2395), .D(R2_n487), .Q(R2_n1391) );
  DLH_X1 R2_shift_in_data_reg_4_ ( .G(R2_n2396), .D(R2_n486), .Q(R2_n1390) );
  DLH_X1 R2_shift_in_data_reg_3_ ( .G(R2_n2395), .D(R2_n485), .Q(R2_n1389) );
  DLH_X1 R2_shift_in_data_reg_2_ ( .G(R2_U22_Z_1), .D(R2_n484), .Q(R2_n1388)
         );
  DLH_X1 R2_shift_in_data_reg_1_ ( .G(R2_n2395), .D(R2_n483), .Q(R2_n1387) );
  DLH_X1 R2_shift_in_data_reg_0_ ( .G(R2_n2396), .D(R2_n482), .Q(R2_n1386) );
  DLH_X1 R2_shift_in_data_reg_99_ ( .G(R2_n2397), .D(R2_n581), .Q(R2_n1485) );
  DLH_X1 R2_shift_in_data_reg_100_ ( .G(R2_U22_Z_1), .D(R2_n582), .Q(R2_n1486)
         );
  DLH_X1 R2_shift_in_data_reg_101_ ( .G(R2_U22_Z_1), .D(R2_n583), .Q(R2_n1487)
         );
  DLH_X1 R2_shift_in_data_reg_102_ ( .G(R2_n2395), .D(R2_n584), .Q(R2_n1488)
         );
  DLH_X1 R2_shift_in_data_reg_103_ ( .G(R2_n2395), .D(R2_n585), .Q(R2_n1489)
         );
  DLH_X1 R2_shift_in_data_reg_104_ ( .G(R2_U22_Z_1), .D(R2_n586), .Q(R2_n1490)
         );
  DLH_X1 R2_shift_in_data_reg_105_ ( .G(R2_n2397), .D(R2_n587), .Q(R2_n1491)
         );
  DLH_X1 R2_shift_in_data_reg_106_ ( .G(R2_n2397), .D(R2_n588), .Q(R2_n1492)
         );
  DLH_X1 R2_shift_in_data_reg_107_ ( .G(R2_n2395), .D(R2_n589), .Q(R2_n1493)
         );
  DLH_X1 R2_shift_in_data_reg_108_ ( .G(R2_n2396), .D(R2_n590), .Q(R2_n1494)
         );
  DLH_X1 R2_shift_in_data_reg_109_ ( .G(R2_n2397), .D(R2_n591), .Q(R2_n1495)
         );
  DLH_X1 R2_shift_in_data_reg_110_ ( .G(R2_n2396), .D(R2_n592), .Q(R2_n1496)
         );
  DLH_X1 R2_shift_in_data_reg_111_ ( .G(R2_n2397), .D(R2_n593), .Q(R2_n1497)
         );
  DLH_X1 R2_shift_in_data_reg_112_ ( .G(R2_n2397), .D(R2_n594), .Q(R2_n1498)
         );
  DLH_X1 R2_shift_in_data_reg_113_ ( .G(R2_n2397), .D(R2_n595), .Q(R2_n1499)
         );
  DLH_X1 R2_shift_in_data_reg_114_ ( .G(R2_n2397), .D(R2_n596), .Q(R2_n1500)
         );
  DLH_X1 R2_shift_in_data_reg_115_ ( .G(R2_n2397), .D(R2_n597), .Q(R2_n1501)
         );
  DLH_X1 R2_shift_in_data_reg_116_ ( .G(R2_n2396), .D(R2_n598), .Q(R2_n1502)
         );
  DLH_X1 R2_shift_in_data_reg_117_ ( .G(R2_n2396), .D(R2_n599), .Q(R2_n1503)
         );
  DLH_X1 R2_shift_in_data_reg_118_ ( .G(R2_n2396), .D(R2_n600), .Q(R2_n1504)
         );
  DLH_X1 R2_shift_in_data_reg_119_ ( .G(R2_n2397), .D(R2_n601), .Q(R2_n1505)
         );
  DLH_X1 R2_shift_in_data_reg_120_ ( .G(R2_n2396), .D(R2_n602), .Q(R2_n1506)
         );
  DLH_X1 R2_shift_in_data_reg_121_ ( .G(R2_n2396), .D(R2_n603), .Q(R2_n1507)
         );
  DLH_X1 R2_shift_in_data_reg_122_ ( .G(R2_n2397), .D(R2_n604), .Q(R2_n1508)
         );
  DLH_X1 R2_shift_in_data_reg_123_ ( .G(R2_n2396), .D(R2_n605), .Q(R2_n1509)
         );
  DLH_X1 R2_shift_in_data_reg_124_ ( .G(R2_n2397), .D(R2_n606), .Q(R2_n1510)
         );
  DLH_X1 R2_shift_in_data_reg_125_ ( .G(R2_n2397), .D(R2_n607), .Q(R2_n1511)
         );
  DLH_X1 R2_shift_in_data_reg_126_ ( .G(R2_n2396), .D(R2_n608), .Q(R2_n1512)
         );
  DLH_X1 R2_shift_in_data_reg_127_ ( .G(R2_n2396), .D(R2_n609), .Q(R2_n1513)
         );
  DFF_X1 R2_temp_sub_data_reg_127_ ( .D(R2_n129), .CK(clk), .Q(R2_n609) );
  DFF_X1 R2_temp_sub_data_reg_126_ ( .D(R2_n128), .CK(clk), .Q(R2_n608) );
  DFF_X1 R2_temp_sub_data_reg_125_ ( .D(R2_n127), .CK(clk), .Q(R2_n607) );
  DFF_X1 R2_temp_sub_data_reg_124_ ( .D(R2_n126), .CK(clk), .Q(R2_n606) );
  DFF_X1 R2_temp_sub_data_reg_123_ ( .D(R2_n125), .CK(clk), .Q(R2_n605) );
  DFF_X1 R2_temp_sub_data_reg_122_ ( .D(R2_n124), .CK(clk), .Q(R2_n604) );
  DFF_X1 R2_temp_sub_data_reg_121_ ( .D(R2_n123), .CK(clk), .Q(R2_n603) );
  DFF_X1 R2_temp_sub_data_reg_120_ ( .D(R2_n122), .CK(clk), .Q(R2_n602) );
  DFF_X1 R2_temp_sub_data_reg_119_ ( .D(R2_n121), .CK(clk), .Q(R2_n601) );
  DFF_X1 R2_temp_sub_data_reg_118_ ( .D(R2_n120), .CK(clk), .Q(R2_n600) );
  DFF_X1 R2_temp_sub_data_reg_117_ ( .D(R2_n119), .CK(clk), .Q(R2_n599) );
  DFF_X1 R2_temp_sub_data_reg_116_ ( .D(R2_n118), .CK(clk), .Q(R2_n598) );
  DFF_X1 R2_temp_sub_data_reg_115_ ( .D(R2_n117), .CK(clk), .Q(R2_n597) );
  DFF_X1 R2_temp_sub_data_reg_114_ ( .D(R2_n116), .CK(clk), .Q(R2_n596) );
  DFF_X1 R2_temp_sub_data_reg_113_ ( .D(R2_n115), .CK(clk), .Q(R2_n595) );
  DFF_X1 R2_temp_sub_data_reg_112_ ( .D(R2_n114), .CK(clk), .Q(R2_n594) );
  DFF_X1 R2_temp_sub_data_reg_111_ ( .D(R2_n113), .CK(clk), .Q(R2_n593) );
  DFF_X1 R2_temp_sub_data_reg_110_ ( .D(R2_n112), .CK(clk), .Q(R2_n592) );
  DFF_X1 R2_temp_sub_data_reg_109_ ( .D(R2_n111), .CK(clk), .Q(R2_n591) );
  DFF_X1 R2_temp_sub_data_reg_108_ ( .D(R2_n110), .CK(clk), .Q(R2_n590) );
  DFF_X1 R2_temp_sub_data_reg_107_ ( .D(R2_n109), .CK(clk), .Q(R2_n589) );
  DFF_X1 R2_temp_sub_data_reg_106_ ( .D(R2_n108), .CK(clk), .Q(R2_n588) );
  DFF_X1 R2_temp_sub_data_reg_105_ ( .D(R2_n107), .CK(clk), .Q(R2_n587) );
  DFF_X1 R2_temp_sub_data_reg_104_ ( .D(R2_n106), .CK(clk), .Q(R2_n586) );
  DFF_X1 R2_temp_sub_data_reg_103_ ( .D(R2_n105), .CK(clk), .Q(R2_n585) );
  DFF_X1 R2_temp_sub_data_reg_102_ ( .D(R2_n104), .CK(clk), .Q(R2_n584) );
  DFF_X1 R2_temp_sub_data_reg_101_ ( .D(R2_n103), .CK(clk), .Q(R2_n583) );
  DFF_X1 R2_temp_sub_data_reg_100_ ( .D(R2_n102), .CK(clk), .Q(R2_n582) );
  DFF_X1 R2_temp_sub_data_reg_99_ ( .D(R2_n101), .CK(clk), .Q(R2_n581) );
  DFF_X1 R2_temp_sub_data_reg_98_ ( .D(R2_n100), .CK(clk), .Q(R2_n580) );
  DFF_X1 R2_temp_sub_data_reg_97_ ( .D(R2_n99), .CK(clk), .Q(R2_n579) );
  DFF_X1 R2_temp_sub_data_reg_96_ ( .D(R2_n98), .CK(clk), .Q(R2_n578) );
  DFF_X1 R2_temp_sub_data_reg_95_ ( .D(R2_n97), .CK(clk), .Q(R2_n577) );
  DFF_X1 R2_temp_sub_data_reg_94_ ( .D(R2_n96), .CK(clk), .Q(R2_n576) );
  DFF_X1 R2_temp_sub_data_reg_93_ ( .D(R2_n95), .CK(clk), .Q(R2_n575) );
  DFF_X1 R2_temp_sub_data_reg_92_ ( .D(R2_n94), .CK(clk), .Q(R2_n574) );
  DFF_X1 R2_temp_sub_data_reg_91_ ( .D(R2_n93), .CK(clk), .Q(R2_n573) );
  DFF_X1 R2_temp_sub_data_reg_90_ ( .D(R2_n92), .CK(clk), .Q(R2_n572) );
  DFF_X1 R2_temp_sub_data_reg_89_ ( .D(R2_n91), .CK(clk), .Q(R2_n571) );
  DFF_X1 R2_temp_sub_data_reg_88_ ( .D(R2_n90), .CK(clk), .Q(R2_n570) );
  DFF_X1 R2_temp_sub_data_reg_87_ ( .D(R2_n89), .CK(clk), .Q(R2_n569) );
  DFF_X1 R2_temp_sub_data_reg_86_ ( .D(R2_n88), .CK(clk), .Q(R2_n568) );
  DFF_X1 R2_temp_sub_data_reg_85_ ( .D(R2_n87), .CK(clk), .Q(R2_n567) );
  DFF_X1 R2_temp_sub_data_reg_84_ ( .D(R2_n86), .CK(clk), .Q(R2_n566) );
  DFF_X1 R2_temp_sub_data_reg_83_ ( .D(R2_n85), .CK(clk), .Q(R2_n565) );
  DFF_X1 R2_temp_sub_data_reg_82_ ( .D(R2_n84), .CK(clk), .Q(R2_n564) );
  DFF_X1 R2_temp_sub_data_reg_81_ ( .D(R2_n83), .CK(clk), .Q(R2_n563) );
  DFF_X1 R2_temp_sub_data_reg_80_ ( .D(R2_n82), .CK(clk), .Q(R2_n562) );
  DFF_X1 R2_temp_sub_data_reg_79_ ( .D(R2_n81), .CK(clk), .Q(R2_n561) );
  DFF_X1 R2_temp_sub_data_reg_78_ ( .D(R2_n80), .CK(clk), .Q(R2_n560) );
  DFF_X1 R2_temp_sub_data_reg_77_ ( .D(R2_n79), .CK(clk), .Q(R2_n559) );
  DFF_X1 R2_temp_sub_data_reg_76_ ( .D(R2_n78), .CK(clk), .Q(R2_n558) );
  DFF_X1 R2_temp_sub_data_reg_75_ ( .D(R2_n77), .CK(clk), .Q(R2_n557) );
  DFF_X1 R2_temp_sub_data_reg_74_ ( .D(R2_n76), .CK(clk), .Q(R2_n556) );
  DFF_X1 R2_temp_sub_data_reg_73_ ( .D(R2_n75), .CK(clk), .Q(R2_n555) );
  DFF_X1 R2_temp_sub_data_reg_72_ ( .D(R2_n74), .CK(clk), .Q(R2_n554) );
  DFF_X1 R2_temp_sub_data_reg_71_ ( .D(R2_n73), .CK(clk), .Q(R2_n553) );
  DFF_X1 R2_temp_sub_data_reg_70_ ( .D(R2_n72), .CK(clk), .Q(R2_n552) );
  DFF_X1 R2_temp_sub_data_reg_69_ ( .D(R2_n71), .CK(clk), .Q(R2_n551) );
  DFF_X1 R2_temp_sub_data_reg_68_ ( .D(R2_n70), .CK(clk), .Q(R2_n550) );
  DFF_X1 R2_temp_sub_data_reg_67_ ( .D(R2_n69), .CK(clk), .Q(R2_n549) );
  DFF_X1 R2_temp_sub_data_reg_66_ ( .D(R2_n68), .CK(clk), .Q(R2_n548) );
  DFF_X1 R2_temp_sub_data_reg_65_ ( .D(R2_n67), .CK(clk), .Q(R2_n547) );
  DFF_X1 R2_temp_sub_data_reg_64_ ( .D(R2_n66), .CK(clk), .Q(R2_n546) );
  DFF_X1 R2_temp_sub_data_reg_63_ ( .D(R2_n65), .CK(clk), .Q(R2_n545) );
  DFF_X1 R2_temp_sub_data_reg_62_ ( .D(R2_n64), .CK(clk), .Q(R2_n544) );
  DFF_X1 R2_temp_sub_data_reg_61_ ( .D(R2_n63), .CK(clk), .Q(R2_n543) );
  DFF_X1 R2_temp_sub_data_reg_60_ ( .D(R2_n62), .CK(clk), .Q(R2_n542) );
  DFF_X1 R2_temp_sub_data_reg_59_ ( .D(R2_n61), .CK(clk), .Q(R2_n541) );
  DFF_X1 R2_temp_sub_data_reg_58_ ( .D(R2_n60), .CK(clk), .Q(R2_n540) );
  DFF_X1 R2_temp_sub_data_reg_57_ ( .D(R2_n59), .CK(clk), .Q(R2_n539) );
  DFF_X1 R2_temp_sub_data_reg_56_ ( .D(R2_n58), .CK(clk), .Q(R2_n538) );
  DFF_X1 R2_temp_sub_data_reg_55_ ( .D(R2_n57), .CK(clk), .Q(R2_n537) );
  DFF_X1 R2_temp_sub_data_reg_54_ ( .D(R2_n56), .CK(clk), .Q(R2_n536) );
  DFF_X1 R2_temp_sub_data_reg_53_ ( .D(R2_n55), .CK(clk), .Q(R2_n535) );
  DFF_X1 R2_temp_sub_data_reg_52_ ( .D(R2_n54), .CK(clk), .Q(R2_n534) );
  DFF_X1 R2_temp_sub_data_reg_51_ ( .D(R2_n53), .CK(clk), .Q(R2_n533) );
  DFF_X1 R2_temp_sub_data_reg_50_ ( .D(R2_n52), .CK(clk), .Q(R2_n532) );
  DFF_X1 R2_temp_sub_data_reg_49_ ( .D(R2_n51), .CK(clk), .Q(R2_n531) );
  DFF_X1 R2_temp_sub_data_reg_48_ ( .D(R2_n50), .CK(clk), .Q(R2_n530) );
  DFF_X1 R2_temp_sub_data_reg_47_ ( .D(R2_n49), .CK(clk), .Q(R2_n529) );
  DFF_X1 R2_temp_sub_data_reg_46_ ( .D(R2_n48), .CK(clk), .Q(R2_n528) );
  DFF_X1 R2_temp_sub_data_reg_45_ ( .D(R2_n47), .CK(clk), .Q(R2_n527) );
  DFF_X1 R2_temp_sub_data_reg_44_ ( .D(R2_n46), .CK(clk), .Q(R2_n526) );
  DFF_X1 R2_temp_sub_data_reg_43_ ( .D(R2_n45), .CK(clk), .Q(R2_n525) );
  DFF_X1 R2_temp_sub_data_reg_42_ ( .D(R2_n44), .CK(clk), .Q(R2_n524) );
  DFF_X1 R2_temp_sub_data_reg_41_ ( .D(R2_n43), .CK(clk), .Q(R2_n523) );
  DFF_X1 R2_temp_sub_data_reg_40_ ( .D(R2_n42), .CK(clk), .Q(R2_n522) );
  DFF_X1 R2_temp_sub_data_reg_39_ ( .D(R2_n41), .CK(clk), .Q(R2_n521) );
  DFF_X1 R2_temp_sub_data_reg_38_ ( .D(R2_n40), .CK(clk), .Q(R2_n520) );
  DFF_X1 R2_temp_sub_data_reg_37_ ( .D(R2_n39), .CK(clk), .Q(R2_n519) );
  DFF_X1 R2_temp_sub_data_reg_36_ ( .D(R2_n38), .CK(clk), .Q(R2_n518) );
  DFF_X1 R2_temp_sub_data_reg_35_ ( .D(R2_n37), .CK(clk), .Q(R2_n517) );
  DFF_X1 R2_temp_sub_data_reg_34_ ( .D(R2_n36), .CK(clk), .Q(R2_n516) );
  DFF_X1 R2_temp_sub_data_reg_33_ ( .D(R2_n35), .CK(clk), .Q(R2_n515) );
  DFF_X1 R2_temp_sub_data_reg_32_ ( .D(R2_n34), .CK(clk), .Q(R2_n514) );
  DFF_X1 R2_temp_sub_data_reg_31_ ( .D(R2_n33), .CK(clk), .Q(R2_n513) );
  DFF_X1 R2_temp_sub_data_reg_30_ ( .D(R2_n32), .CK(clk), .Q(R2_n512) );
  DFF_X1 R2_temp_sub_data_reg_29_ ( .D(R2_n31), .CK(clk), .Q(R2_n511) );
  DFF_X1 R2_temp_sub_data_reg_28_ ( .D(R2_n30), .CK(clk), .Q(R2_n510) );
  DFF_X1 R2_temp_sub_data_reg_27_ ( .D(R2_n29), .CK(clk), .Q(R2_n509) );
  DFF_X1 R2_temp_sub_data_reg_26_ ( .D(R2_n28), .CK(clk), .Q(R2_n508) );
  DFF_X1 R2_temp_sub_data_reg_25_ ( .D(R2_n27), .CK(clk), .Q(R2_n507) );
  DFF_X1 R2_temp_sub_data_reg_24_ ( .D(R2_n26), .CK(clk), .Q(R2_n506) );
  DFF_X1 R2_temp_sub_data_reg_23_ ( .D(R2_n25), .CK(clk), .Q(R2_n505) );
  DFF_X1 R2_temp_sub_data_reg_22_ ( .D(R2_n24), .CK(clk), .Q(R2_n504) );
  DFF_X1 R2_temp_sub_data_reg_21_ ( .D(R2_n23), .CK(clk), .Q(R2_n503) );
  DFF_X1 R2_temp_sub_data_reg_20_ ( .D(R2_n22), .CK(clk), .Q(R2_n502) );
  DFF_X1 R2_temp_sub_data_reg_19_ ( .D(R2_n21), .CK(clk), .Q(R2_n501) );
  DFF_X1 R2_temp_sub_data_reg_18_ ( .D(R2_n20), .CK(clk), .Q(R2_n500) );
  DFF_X1 R2_temp_sub_data_reg_17_ ( .D(R2_n19), .CK(clk), .Q(R2_n499) );
  DFF_X1 R2_temp_sub_data_reg_16_ ( .D(R2_n18), .CK(clk), .Q(R2_n498) );
  DFF_X1 R2_temp_sub_data_reg_15_ ( .D(R2_n17), .CK(clk), .Q(R2_n497) );
  DFF_X1 R2_temp_sub_data_reg_14_ ( .D(R2_n16), .CK(clk), .Q(R2_n496) );
  DFF_X1 R2_temp_sub_data_reg_13_ ( .D(R2_n15), .CK(clk), .Q(R2_n495) );
  DFF_X1 R2_temp_sub_data_reg_12_ ( .D(R2_n14), .CK(clk), .Q(R2_n494) );
  DFF_X1 R2_temp_sub_data_reg_11_ ( .D(R2_n13), .CK(clk), .Q(R2_n493) );
  DFF_X1 R2_temp_sub_data_reg_10_ ( .D(R2_n12), .CK(clk), .Q(R2_n492) );
  DFF_X1 R2_temp_sub_data_reg_9_ ( .D(R2_n11), .CK(clk), .Q(R2_n491) );
  DFF_X1 R2_temp_sub_data_reg_8_ ( .D(R2_n10), .CK(clk), .Q(R2_n490) );
  DFF_X1 R2_temp_sub_data_reg_7_ ( .D(R2_n9), .CK(clk), .Q(R2_n489) );
  DFF_X1 R2_temp_sub_data_reg_6_ ( .D(R2_n8), .CK(clk), .Q(R2_n488) );
  DFF_X1 R2_temp_sub_data_reg_5_ ( .D(R2_n7), .CK(clk), .Q(R2_n487) );
  DFF_X1 R2_temp_sub_data_reg_4_ ( .D(R2_n6), .CK(clk), .Q(R2_n486) );
  DFF_X1 R2_temp_sub_data_reg_3_ ( .D(R2_n5), .CK(clk), .Q(R2_n485) );
  DFF_X1 R2_temp_sub_data_reg_2_ ( .D(R2_n4), .CK(clk), .Q(R2_n484) );
  DFF_X1 R2_temp_sub_data_reg_1_ ( .D(R2_n3), .CK(clk), .Q(R2_n483) );
  DFF_X1 R2_temp_sub_data_reg_0_ ( .D(R2_n2), .CK(clk), .Q(R2_n482) );
  DFF_X1 R2_cnt_reg_3_ ( .D(R2_n2341), .CK(clk), .Q(R2_r332_A_3_) );
  DFF_X1 R2_cnt_reg_2_ ( .D(R2_n2340), .CK(clk), .Q(R2_r332_A_2_), .QN(
        R2_n1804) );
  DFF_X1 R2_cnt_reg_1_ ( .D(R2_n2339), .CK(clk), .Q(R2_r332_A_1_), .QN(
        R2_n1805) );
  DFF_X1 R2_cnt_reg_0_ ( .D(R2_n2338), .CK(clk), .Q(R2_r332_A_0_), .QN(
        R2_n1806) );
  DLH_X1 R2_sub_in_data_reg_98_ ( .G(R2_n2405), .D(n3618), .Q(R2_n1742) );
  DLH_X1 R2_sub_in_data_reg_97_ ( .G(R2_n2407), .D(n3617), .Q(R2_n1741) );
  DLH_X1 R2_sub_in_data_reg_96_ ( .G(R2_n2405), .D(n3616), .Q(R2_n1740) );
  DLH_X1 R2_sub_in_data_reg_95_ ( .G(R2_n2406), .D(n3615), .Q(R2_n1739) );
  DLH_X1 R2_sub_in_data_reg_94_ ( .G(R2_U24_Z_1), .D(n3614), .Q(R2_n1738) );
  DLH_X1 R2_sub_in_data_reg_93_ ( .G(R2_U24_Z_1), .D(n3613), .Q(R2_n1737) );
  DLH_X1 R2_sub_in_data_reg_92_ ( .G(R2_n2406), .D(n3612), .Q(R2_n1736) );
  DLH_X1 R2_sub_in_data_reg_91_ ( .G(R2_n2405), .D(n3611), .Q(R2_n1735) );
  DLH_X1 R2_sub_in_data_reg_90_ ( .G(R2_U24_Z_1), .D(n3610), .Q(R2_n1734) );
  DLH_X1 R2_sub_in_data_reg_89_ ( .G(R2_U24_Z_1), .D(n3609), .Q(R2_n1733) );
  DLH_X1 R2_sub_in_data_reg_88_ ( .G(R2_U24_Z_1), .D(n3608), .Q(R2_n1732) );
  DLH_X1 R2_sub_in_data_reg_87_ ( .G(R2_n2407), .D(n3607), .Q(R2_n1731) );
  DLH_X1 R2_sub_in_data_reg_86_ ( .G(R2_U24_Z_1), .D(n3606), .Q(R2_n1730) );
  DLH_X1 R2_sub_in_data_reg_85_ ( .G(R2_n2406), .D(n3605), .Q(R2_n1729) );
  DLH_X1 R2_sub_in_data_reg_84_ ( .G(R2_U24_Z_1), .D(n3604), .Q(R2_n1728) );
  DLH_X1 R2_sub_in_data_reg_83_ ( .G(R2_n2405), .D(n3603), .Q(R2_n1727) );
  DLH_X1 R2_sub_in_data_reg_82_ ( .G(R2_n2407), .D(n3602), .Q(R2_n1726) );
  DLH_X1 R2_sub_in_data_reg_81_ ( .G(R2_n2406), .D(n3601), .Q(R2_n1725) );
  DLH_X1 R2_sub_in_data_reg_80_ ( .G(R2_n2405), .D(n3600), .Q(R2_n1724) );
  DLH_X1 R2_sub_in_data_reg_79_ ( .G(R2_n2405), .D(n3599), .Q(R2_n1723) );
  DLH_X1 R2_sub_in_data_reg_78_ ( .G(R2_n2405), .D(n3598), .Q(R2_n1722) );
  DLH_X1 R2_sub_in_data_reg_77_ ( .G(R2_n2405), .D(n3597), .Q(R2_n1721) );
  DLH_X1 R2_sub_in_data_reg_76_ ( .G(R2_U24_Z_1), .D(n3596), .Q(R2_n1720) );
  DLH_X1 R2_sub_in_data_reg_75_ ( .G(R2_n2407), .D(n3595), .Q(R2_n1719) );
  DLH_X1 R2_sub_in_data_reg_74_ ( .G(R2_U24_Z_1), .D(n3594), .Q(R2_n1718) );
  DLH_X1 R2_sub_in_data_reg_73_ ( .G(R2_n2407), .D(n3593), .Q(R2_n1717) );
  DLH_X1 R2_sub_in_data_reg_72_ ( .G(R2_n2407), .D(n3592), .Q(R2_n1716) );
  DLH_X1 R2_sub_in_data_reg_71_ ( .G(R2_n2406), .D(n3591), .Q(R2_n1715) );
  DLH_X1 R2_sub_in_data_reg_70_ ( .G(R2_n2406), .D(n3590), .Q(R2_n1714) );
  DLH_X1 R2_sub_in_data_reg_69_ ( .G(R2_n2405), .D(n3589), .Q(R2_n1713) );
  DLH_X1 R2_sub_in_data_reg_68_ ( .G(R2_n2406), .D(n3588), .Q(R2_n1712) );
  DLH_X1 R2_sub_in_data_reg_67_ ( .G(R2_n2406), .D(n3587), .Q(R2_n1711) );
  DLH_X1 R2_sub_in_data_reg_66_ ( .G(R2_n2407), .D(n3586), .Q(R2_n1710) );
  DLH_X1 R2_sub_in_data_reg_65_ ( .G(R2_n2405), .D(n3585), .Q(R2_n1709) );
  DLH_X1 R2_sub_in_data_reg_64_ ( .G(R2_U24_Z_1), .D(n3584), .Q(R2_n1708) );
  DLH_X1 R2_sub_in_data_reg_63_ ( .G(R2_n2405), .D(n3583), .Q(R2_n1707) );
  DLH_X1 R2_sub_in_data_reg_62_ ( .G(R2_n2406), .D(n3582), .Q(R2_n1706) );
  DLH_X1 R2_sub_in_data_reg_61_ ( .G(R2_U24_Z_1), .D(n3581), .Q(R2_n1705) );
  DLH_X1 R2_sub_in_data_reg_60_ ( .G(R2_n2406), .D(n3580), .Q(R2_n1704) );
  DLH_X1 R2_sub_in_data_reg_59_ ( .G(R2_n2407), .D(n3579), .Q(R2_n1703) );
  DLH_X1 R2_sub_in_data_reg_58_ ( .G(R2_n2406), .D(n3578), .Q(R2_n1702) );
  DLH_X1 R2_sub_in_data_reg_57_ ( .G(R2_n2407), .D(n3577), .Q(R2_n1701) );
  DLH_X1 R2_sub_in_data_reg_56_ ( .G(R2_n2407), .D(n3576), .Q(R2_n1700) );
  DLH_X1 R2_sub_in_data_reg_55_ ( .G(R2_n2406), .D(n3575), .Q(R2_n1699) );
  DLH_X1 R2_sub_in_data_reg_54_ ( .G(R2_n2405), .D(n3574), .Q(R2_n1698) );
  DLH_X1 R2_sub_in_data_reg_53_ ( .G(R2_U24_Z_1), .D(n3573), .Q(R2_n1697) );
  DLH_X1 R2_sub_in_data_reg_52_ ( .G(R2_n2405), .D(n3572), .Q(R2_n1696) );
  DLH_X1 R2_sub_in_data_reg_51_ ( .G(R2_U24_Z_1), .D(n3571), .Q(R2_n1695) );
  DLH_X1 R2_sub_in_data_reg_50_ ( .G(R2_U24_Z_1), .D(n3570), .Q(R2_n1694) );
  DLH_X1 R2_sub_in_data_reg_49_ ( .G(R2_n2407), .D(n3569), .Q(R2_n1693) );
  DLH_X1 R2_sub_in_data_reg_48_ ( .G(R2_n2405), .D(n3568), .Q(R2_n1692) );
  DLH_X1 R2_sub_in_data_reg_47_ ( .G(R2_U24_Z_1), .D(n3567), .Q(R2_n1691) );
  DLH_X1 R2_sub_in_data_reg_46_ ( .G(R2_n2407), .D(n3566), .Q(R2_n1690) );
  DLH_X1 R2_sub_in_data_reg_45_ ( .G(R2_n2406), .D(n3565), .Q(R2_n1689) );
  DLH_X1 R2_sub_in_data_reg_44_ ( .G(R2_n2407), .D(n3564), .Q(R2_n1688) );
  DLH_X1 R2_sub_in_data_reg_43_ ( .G(R2_U24_Z_1), .D(n3563), .Q(R2_n1687) );
  DLH_X1 R2_sub_in_data_reg_42_ ( .G(R2_U24_Z_1), .D(n3562), .Q(R2_n1686) );
  DLH_X1 R2_sub_in_data_reg_41_ ( .G(R2_n2407), .D(n3561), .Q(R2_n1685) );
  DLH_X1 R2_sub_in_data_reg_40_ ( .G(R2_U24_Z_1), .D(n3560), .Q(R2_n1684) );
  DLH_X1 R2_sub_in_data_reg_39_ ( .G(R2_n2407), .D(n3559), .Q(R2_n1683) );
  DLH_X1 R2_sub_in_data_reg_38_ ( .G(R2_n2406), .D(n3558), .Q(R2_n1682) );
  DLH_X1 R2_sub_in_data_reg_37_ ( .G(R2_n2406), .D(n3557), .Q(R2_n1681) );
  DLH_X1 R2_sub_in_data_reg_36_ ( .G(R2_n2405), .D(n3556), .Q(R2_n1680) );
  DLH_X1 R2_sub_in_data_reg_35_ ( .G(R2_n2405), .D(n3555), .Q(R2_n1679) );
  DLH_X1 R2_sub_in_data_reg_34_ ( .G(R2_n2405), .D(n3554), .Q(R2_n1678) );
  DLH_X1 R2_sub_in_data_reg_33_ ( .G(R2_U24_Z_1), .D(n3553), .Q(R2_n1677) );
  DLH_X1 R2_sub_in_data_reg_32_ ( .G(R2_n2405), .D(n3552), .Q(R2_n1676) );
  DLH_X1 R2_sub_in_data_reg_31_ ( .G(R2_n2405), .D(n3551), .Q(R2_n1675) );
  DLH_X1 R2_sub_in_data_reg_30_ ( .G(R2_n2405), .D(n3550), .Q(R2_n1674) );
  DLH_X1 R2_sub_in_data_reg_29_ ( .G(R2_n2405), .D(n3549), .Q(R2_n1673) );
  DLH_X1 R2_sub_in_data_reg_28_ ( .G(R2_n2405), .D(n3548), .Q(R2_n1672) );
  DLH_X1 R2_sub_in_data_reg_27_ ( .G(R2_n2405), .D(n3547), .Q(R2_n1671) );
  DLH_X1 R2_sub_in_data_reg_26_ ( .G(R2_n2405), .D(n3546), .Q(R2_n1670) );
  DLH_X1 R2_sub_in_data_reg_25_ ( .G(R2_n2405), .D(n3545), .Q(R2_n1669) );
  DLH_X1 R2_sub_in_data_reg_24_ ( .G(R2_n2405), .D(n3544), .Q(R2_n1668) );
  DLH_X1 R2_sub_in_data_reg_23_ ( .G(R2_n2405), .D(n3543), .Q(R2_n1667) );
  DLH_X1 R2_sub_in_data_reg_22_ ( .G(R2_n2405), .D(n3542), .Q(R2_n1666) );
  DLH_X1 R2_sub_in_data_reg_21_ ( .G(R2_n2406), .D(n3541), .Q(R2_n1665) );
  DLH_X1 R2_sub_in_data_reg_20_ ( .G(R2_U24_Z_1), .D(n3540), .Q(R2_n1664) );
  DLH_X1 R2_sub_in_data_reg_19_ ( .G(R2_U24_Z_1), .D(n3539), .Q(R2_n1663) );
  DLH_X1 R2_sub_in_data_reg_18_ ( .G(R2_n2407), .D(n3538), .Q(R2_n1662) );
  DLH_X1 R2_sub_in_data_reg_17_ ( .G(R2_n2406), .D(n3537), .Q(R2_n1661) );
  DLH_X1 R2_sub_in_data_reg_16_ ( .G(R2_U24_Z_1), .D(n3536), .Q(R2_n1660) );
  DLH_X1 R2_sub_in_data_reg_15_ ( .G(R2_n2407), .D(n3535), .Q(R2_n1659) );
  DLH_X1 R2_sub_in_data_reg_14_ ( .G(R2_n2405), .D(n3534), .Q(R2_n1658) );
  DLH_X1 R2_sub_in_data_reg_13_ ( .G(R2_n2407), .D(n3533), .Q(R2_n1657) );
  DLH_X1 R2_sub_in_data_reg_12_ ( .G(R2_n2406), .D(n3532), .Q(R2_n1656) );
  DLH_X1 R2_sub_in_data_reg_11_ ( .G(R2_n2407), .D(n3531), .Q(R2_n1655) );
  DLH_X1 R2_sub_in_data_reg_10_ ( .G(R2_n2406), .D(n3530), .Q(R2_n1654) );
  DLH_X1 R2_sub_in_data_reg_9_ ( .G(R2_n2406), .D(n3529), .Q(R2_n1653) );
  DLH_X1 R2_sub_in_data_reg_8_ ( .G(R2_n2406), .D(n3528), .Q(R2_n1652) );
  DLH_X1 R2_sub_in_data_reg_7_ ( .G(R2_n2406), .D(n3527), .Q(R2_n1651) );
  DLH_X1 R2_sub_in_data_reg_6_ ( .G(R2_n2406), .D(n3526), .Q(R2_n1650) );
  DLH_X1 R2_sub_in_data_reg_5_ ( .G(R2_n2406), .D(n3525), .Q(R2_n1649) );
  DLH_X1 R2_sub_in_data_reg_4_ ( .G(R2_n2406), .D(n3524), .Q(R2_n1648) );
  DLH_X1 R2_sub_in_data_reg_3_ ( .G(R2_n2406), .D(n3523), .Q(R2_n1647) );
  DLH_X1 R2_sub_in_data_reg_2_ ( .G(R2_n2406), .D(n3522), .Q(R2_n1646) );
  DLH_X1 R2_sub_in_data_reg_1_ ( .G(R2_n2406), .D(n3521), .Q(R2_n1645) );
  DLH_X1 R2_sub_in_data_reg_0_ ( .G(R2_n2406), .D(n3520), .Q(R2_n1644) );
  DLH_X1 R2_sub_in_data_reg_99_ ( .G(R2_n2405), .D(n3619), .Q(R2_n1743) );
  DLH_X1 R2_sub_in_data_reg_100_ ( .G(R2_n2407), .D(n3620), .Q(R2_n1744) );
  DLH_X1 R2_sub_in_data_reg_101_ ( .G(R2_n2407), .D(n3621), .Q(R2_n1745) );
  DLH_X1 R2_sub_in_data_reg_102_ ( .G(R2_n2406), .D(n3622), .Q(R2_n1746) );
  DLH_X1 R2_sub_in_data_reg_103_ ( .G(R2_n2406), .D(n3623), .Q(R2_n1747) );
  DLH_X1 R2_sub_in_data_reg_104_ ( .G(R2_n2406), .D(n3624), .Q(R2_n1748) );
  DLH_X1 R2_sub_in_data_reg_105_ ( .G(R2_U24_Z_1), .D(n3625), .Q(R2_n1749) );
  DLH_X1 R2_sub_in_data_reg_106_ ( .G(R2_n2407), .D(n3626), .Q(R2_n1750) );
  DLH_X1 R2_sub_in_data_reg_107_ ( .G(R2_n2405), .D(n3627), .Q(R2_n1751) );
  DLH_X1 R2_sub_in_data_reg_108_ ( .G(R2_n2405), .D(n3628), .Q(R2_n1752) );
  DLH_X1 R2_sub_in_data_reg_109_ ( .G(R2_U24_Z_1), .D(n3629), .Q(R2_n1753) );
  DLH_X1 R2_sub_in_data_reg_110_ ( .G(R2_n2407), .D(n3630), .Q(R2_n1754) );
  DLH_X1 R2_sub_in_data_reg_111_ ( .G(R2_n2407), .D(n3631), .Q(R2_n1755) );
  DLH_X1 R2_sub_in_data_reg_112_ ( .G(R2_n2407), .D(n3632), .Q(R2_n1756) );
  DLH_X1 R2_sub_in_data_reg_113_ ( .G(R2_n2407), .D(n3633), .Q(R2_n1757) );
  DLH_X1 R2_sub_in_data_reg_114_ ( .G(R2_n2407), .D(n3634), .Q(R2_n1758) );
  DLH_X1 R2_sub_in_data_reg_115_ ( .G(R2_n2407), .D(n3635), .Q(R2_n1759) );
  DLH_X1 R2_sub_in_data_reg_116_ ( .G(R2_n2407), .D(n3636), .Q(R2_n1760) );
  DLH_X1 R2_sub_in_data_reg_117_ ( .G(R2_n2407), .D(n3637), .Q(R2_n1761) );
  DLH_X1 R2_sub_in_data_reg_118_ ( .G(R2_n2407), .D(n3638), .Q(R2_n1762) );
  DLH_X1 R2_sub_in_data_reg_119_ ( .G(R2_n2407), .D(n3639), .Q(R2_n1763) );
  DLH_X1 R2_sub_in_data_reg_120_ ( .G(R2_n2407), .D(n3640), .Q(R2_n1764) );
  DLH_X1 R2_sub_in_data_reg_121_ ( .G(R2_U24_Z_1), .D(n3641), .Q(R2_n1765) );
  DLH_X1 R2_sub_in_data_reg_122_ ( .G(R2_U24_Z_1), .D(n3642), .Q(R2_n1766) );
  DLH_X1 R2_sub_in_data_reg_123_ ( .G(R2_U24_Z_1), .D(n3643), .Q(R2_n1767) );
  DLH_X1 R2_sub_in_data_reg_124_ ( .G(R2_U24_Z_1), .D(n3644), .Q(R2_n1768) );
  DLH_X1 R2_sub_in_data_reg_125_ ( .G(R2_U24_Z_1), .D(n3645), .Q(R2_n1769) );
  DLH_X1 R2_sub_in_data_reg_126_ ( .G(R2_U24_Z_1), .D(n3646), .Q(R2_n1770) );
  DLH_X1 R2_sub_in_data_reg_127_ ( .G(R2_U24_Z_1), .D(n3647), .Q(R2_n1771) );
  DLL_X1 R2_temp_round_reg ( .D(n3391), .GN(n3262), .Q(R2_n610) );
  DFF_X1 R2_ready_reg ( .D(R2_n2342), .CK(clk), .Q(n3262), .QN(R2_n1807) );
  SDFF_X1 R2_rstSB_reg ( .D(n3261), .SI(R2_n2346), .SE(R2_n2334), .CK(clk), 
        .Q(R2_n1514) );
  NAND2_X2 R2_SB_U65 ( .A1(R2_SB_n617), .A2(R2_SB_n38), .ZN(R2_SB_n41) );
  CLKBUF_X2 R2_SB_U64 ( .A(R2_SB_n41), .Z(R2_SB_n623) );
  CLKBUF_X2 R2_SB_U60 ( .A(R2_SB_n276), .Z(R2_SB_n628) );
  CLKBUF_X2 R2_SB_U25 ( .A(R2_SB_n628), .Z(R2_SB_n627) );
  AND2_X2 R2_SB_U24 ( .A1(R2_SB_add_108_A_0_), .A2(R2_SB_n442), .ZN(R2_SB_n361) );
  NAND2_X2 R2_SB_U23 ( .A1(R2_SB_n616), .A2(R2_SB_n38), .ZN(R2_SB_n45) );
  CLKBUF_X2 R2_SB_U22 ( .A(R2_SB_n45), .Z(R2_SB_n619) );
  NAND2_X2 R2_SB_U19 ( .A1(R2_SB_n618), .A2(R2_SB_n38), .ZN(R2_SB_n39) );
  CLKBUF_X2 R2_SB_U17 ( .A(R2_SB_n276), .Z(R2_SB_n629) );
  AND2_X2 R2_SB_U10 ( .A1(R2_SB_n442), .A2(R2_SB_n37), .ZN(R2_SB_n363) );
  NOR2_X2 R2_SB_U8 ( .A1(R2_SB_n34), .A2(R2_SB_n37), .ZN(R2_SB_n367) );
  CLKBUF_X2 R2_SB_U5 ( .A(R2_SB_n367), .Z(R2_SB_n616) );
  NAND2_X2 R2_SB_U4 ( .A1(R2_SB_U4_Z_0), .A2(R2_SB_n365), .ZN(R2_SB_n43) );
  NAND2_X2 R2_SB_U3 ( .A1(R2_SB_n615), .A2(R2_SB_n34), .ZN(R2_SB_U11_Z_0) );
  DLH_X2 R2_SB_sbox_s1_reg_1_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_1), .Q(
        R2_SB_n338) );
  DLH_X2 R2_SB_sbox_s2_reg_1_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_1), .Q(
        R2_SB_n322) );
  DLH_X2 R2_SB_sbox_s3_reg_1_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_1), .Q(
        R2_SB_n306) );
  DLH_X2 R2_SB_sbox_s4_reg_1_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_1), .Q(
        R2_SB_n290) );
  DFF_X2 R2_SB_flag_reg ( .D(R2_SB_n571), .CK(clk), .Q(R2_SB_n276) );
  AOI22_X1 R2_SB_U430 ( .A1(R2_n1732), .A2(R2_SB_n363), .B1(R2_n1700), .B2(
        R2_SB_n367), .ZN(R2_SB_n419) );
  AOI22_X1 R2_SB_U429 ( .A1(R2_n1668), .A2(R2_SB_n614), .B1(R2_n1764), .B2(
        R2_SB_n361), .ZN(R2_SB_n418) );
  NAND2_X1 R2_SB_U428 ( .A1(R2_SB_n418), .A2(R2_SB_n419), .ZN(R2_SB_U7_Z_0) );
  AOI22_X1 R2_SB_U427 ( .A1(R2_n1715), .A2(R2_SB_n617), .B1(R2_n1683), .B2(
        R2_SB_n367), .ZN(R2_SB_n427) );
  AOI22_X1 R2_SB_U426 ( .A1(R2_n1651), .A2(R2_SB_n615), .B1(R2_n1747), .B2(
        R2_SB_n618), .ZN(R2_SB_n426) );
  NAND2_X1 R2_SB_U425 ( .A1(R2_SB_n426), .A2(R2_SB_n427), .ZN(R2_SB_U10_Z_7)
         );
  AOI22_X1 R2_SB_U424 ( .A1(R2_n1714), .A2(R2_SB_n617), .B1(R2_n1682), .B2(
        R2_SB_n367), .ZN(R2_SB_n429) );
  AOI22_X1 R2_SB_U423 ( .A1(R2_n1650), .A2(R2_SB_n614), .B1(R2_n1746), .B2(
        R2_SB_n618), .ZN(R2_SB_n428) );
  NAND2_X1 R2_SB_U422 ( .A1(R2_SB_n428), .A2(R2_SB_n429), .ZN(R2_SB_U10_Z_6)
         );
  AOI22_X1 R2_SB_U421 ( .A1(R2_n1713), .A2(R2_SB_n617), .B1(R2_n1681), .B2(
        R2_SB_n367), .ZN(R2_SB_n431) );
  AOI22_X1 R2_SB_U420 ( .A1(R2_n1649), .A2(R2_SB_n373), .B1(R2_n1745), .B2(
        R2_SB_n618), .ZN(R2_SB_n430) );
  NAND2_X1 R2_SB_U419 ( .A1(R2_SB_n430), .A2(R2_SB_n431), .ZN(R2_SB_U10_Z_5)
         );
  AOI22_X1 R2_SB_U418 ( .A1(R2_n1712), .A2(R2_SB_n617), .B1(R2_n1680), .B2(
        R2_SB_n367), .ZN(R2_SB_n433) );
  AOI22_X1 R2_SB_U417 ( .A1(R2_n1648), .A2(R2_SB_n373), .B1(R2_n1744), .B2(
        R2_SB_n618), .ZN(R2_SB_n432) );
  NAND2_X1 R2_SB_U416 ( .A1(R2_SB_n432), .A2(R2_SB_n433), .ZN(R2_SB_U10_Z_4)
         );
  AOI22_X1 R2_SB_U415 ( .A1(R2_n1711), .A2(R2_SB_n617), .B1(R2_n1679), .B2(
        R2_SB_n367), .ZN(R2_SB_n435) );
  AOI22_X1 R2_SB_U413 ( .A1(R2_n1647), .A2(R2_SB_n373), .B1(R2_n1743), .B2(
        R2_SB_n618), .ZN(R2_SB_n434) );
  NAND2_X1 R2_SB_U412 ( .A1(R2_SB_n434), .A2(R2_SB_n435), .ZN(R2_SB_U10_Z_3)
         );
  AOI22_X1 R2_SB_U411 ( .A1(R2_n1710), .A2(R2_SB_n617), .B1(R2_n1678), .B2(
        R2_SB_n367), .ZN(R2_SB_n437) );
  AOI22_X1 R2_SB_U410 ( .A1(R2_n1646), .A2(R2_SB_n373), .B1(R2_n1742), .B2(
        R2_SB_n618), .ZN(R2_SB_n436) );
  NAND2_X1 R2_SB_U409 ( .A1(R2_SB_n436), .A2(R2_SB_n437), .ZN(R2_SB_U10_Z_2)
         );
  AOI22_X1 R2_SB_U408 ( .A1(R2_n1709), .A2(R2_SB_n617), .B1(R2_n1677), .B2(
        R2_SB_n367), .ZN(R2_SB_n439) );
  AOI22_X1 R2_SB_U407 ( .A1(R2_n1645), .A2(R2_SB_n373), .B1(R2_n1741), .B2(
        R2_SB_n618), .ZN(R2_SB_n438) );
  NAND2_X1 R2_SB_U406 ( .A1(R2_SB_n438), .A2(R2_SB_n439), .ZN(R2_SB_U10_Z_1)
         );
  AOI22_X1 R2_SB_U405 ( .A1(R2_n1739), .A2(R2_SB_n363), .B1(R2_n1707), .B2(
        R2_SB_n616), .ZN(R2_SB_n405) );
  AOI22_X1 R2_SB_U404 ( .A1(R2_n1675), .A2(R2_SB_n615), .B1(R2_n1771), .B2(
        R2_SB_n361), .ZN(R2_SB_n404) );
  NAND2_X1 R2_SB_U403 ( .A1(R2_SB_n404), .A2(R2_SB_n405), .ZN(R2_SB_U7_Z_7) );
  AOI22_X1 R2_SB_U402 ( .A1(R2_n1738), .A2(R2_SB_n363), .B1(R2_n1706), .B2(
        R2_SB_n616), .ZN(R2_SB_n407) );
  AOI22_X1 R2_SB_U401 ( .A1(R2_n1674), .A2(R2_SB_n615), .B1(R2_n1770), .B2(
        R2_SB_n361), .ZN(R2_SB_n406) );
  NAND2_X1 R2_SB_U400 ( .A1(R2_SB_n406), .A2(R2_SB_n407), .ZN(R2_SB_U7_Z_6) );
  AOI22_X1 R2_SB_U399 ( .A1(R2_n1737), .A2(R2_SB_n363), .B1(R2_n1705), .B2(
        R2_SB_n616), .ZN(R2_SB_n409) );
  AOI22_X1 R2_SB_U398 ( .A1(R2_n1673), .A2(R2_SB_n615), .B1(R2_n1769), .B2(
        R2_SB_n361), .ZN(R2_SB_n408) );
  NAND2_X1 R2_SB_U397 ( .A1(R2_SB_n408), .A2(R2_SB_n409), .ZN(R2_SB_U7_Z_5) );
  AOI22_X1 R2_SB_U396 ( .A1(R2_n1736), .A2(R2_SB_n363), .B1(R2_n1704), .B2(
        R2_SB_n616), .ZN(R2_SB_n411) );
  AOI22_X1 R2_SB_U395 ( .A1(R2_n1672), .A2(R2_SB_n615), .B1(R2_n1768), .B2(
        R2_SB_n361), .ZN(R2_SB_n410) );
  NAND2_X1 R2_SB_U394 ( .A1(R2_SB_n410), .A2(R2_SB_n411), .ZN(R2_SB_U7_Z_4) );
  AOI22_X1 R2_SB_U393 ( .A1(R2_n1735), .A2(R2_SB_n363), .B1(R2_n1703), .B2(
        R2_SB_n616), .ZN(R2_SB_n413) );
  AOI22_X1 R2_SB_U392 ( .A1(R2_n1671), .A2(R2_SB_n615), .B1(R2_n1767), .B2(
        R2_SB_n361), .ZN(R2_SB_n412) );
  NAND2_X1 R2_SB_U391 ( .A1(R2_SB_n412), .A2(R2_SB_n413), .ZN(R2_SB_U7_Z_3) );
  AOI22_X1 R2_SB_U390 ( .A1(R2_n1734), .A2(R2_SB_n363), .B1(R2_n1702), .B2(
        R2_SB_n367), .ZN(R2_SB_n415) );
  AOI22_X1 R2_SB_U389 ( .A1(R2_n1670), .A2(R2_SB_n615), .B1(R2_n1766), .B2(
        R2_SB_n361), .ZN(R2_SB_n414) );
  NAND2_X1 R2_SB_U388 ( .A1(R2_SB_n414), .A2(R2_SB_n415), .ZN(R2_SB_U7_Z_2) );
  AOI22_X1 R2_SB_U387 ( .A1(R2_n1733), .A2(R2_SB_n363), .B1(R2_n1701), .B2(
        R2_SB_n367), .ZN(R2_SB_n417) );
  AOI22_X1 R2_SB_U386 ( .A1(R2_n1669), .A2(R2_SB_n615), .B1(R2_n1765), .B2(
        R2_SB_n361), .ZN(R2_SB_n416) );
  NAND2_X1 R2_SB_U385 ( .A1(R2_SB_n416), .A2(R2_SB_n417), .ZN(R2_SB_U7_Z_1) );
  AOI22_X1 R2_SB_U384 ( .A1(R2_n1731), .A2(R2_SB_n363), .B1(R2_n1699), .B2(
        R2_SB_n616), .ZN(R2_SB_n389) );
  AOI22_X1 R2_SB_U383 ( .A1(R2_n1667), .A2(R2_SB_n614), .B1(R2_n1763), .B2(
        R2_SB_n361), .ZN(R2_SB_n388) );
  NAND2_X1 R2_SB_U382 ( .A1(R2_SB_n388), .A2(R2_SB_n389), .ZN(R2_SB_U8_Z_7) );
  AOI22_X1 R2_SB_U381 ( .A1(R2_n1730), .A2(R2_SB_n363), .B1(R2_n1698), .B2(
        R2_SB_n616), .ZN(R2_SB_n391) );
  AOI22_X1 R2_SB_U380 ( .A1(R2_n1666), .A2(R2_SB_n614), .B1(R2_n1762), .B2(
        R2_SB_n361), .ZN(R2_SB_n390) );
  NAND2_X1 R2_SB_U379 ( .A1(R2_SB_n390), .A2(R2_SB_n391), .ZN(R2_SB_U8_Z_6) );
  AOI22_X1 R2_SB_U378 ( .A1(R2_n1729), .A2(R2_SB_n363), .B1(R2_n1697), .B2(
        R2_SB_n616), .ZN(R2_SB_n393) );
  AOI22_X1 R2_SB_U377 ( .A1(R2_n1665), .A2(R2_SB_n614), .B1(R2_n1761), .B2(
        R2_SB_n361), .ZN(R2_SB_n392) );
  NAND2_X1 R2_SB_U376 ( .A1(R2_SB_n392), .A2(R2_SB_n393), .ZN(R2_SB_U8_Z_5) );
  AOI22_X1 R2_SB_U375 ( .A1(R2_n1728), .A2(R2_SB_n363), .B1(R2_n1696), .B2(
        R2_SB_n616), .ZN(R2_SB_n395) );
  AOI22_X1 R2_SB_U374 ( .A1(R2_n1664), .A2(R2_SB_n614), .B1(R2_n1760), .B2(
        R2_SB_n361), .ZN(R2_SB_n394) );
  NAND2_X1 R2_SB_U373 ( .A1(R2_SB_n394), .A2(R2_SB_n395), .ZN(R2_SB_U8_Z_4) );
  AOI22_X1 R2_SB_U372 ( .A1(R2_n1727), .A2(R2_SB_n363), .B1(R2_n1695), .B2(
        R2_SB_n616), .ZN(R2_SB_n397) );
  AOI22_X1 R2_SB_U371 ( .A1(R2_n1663), .A2(R2_SB_n615), .B1(R2_n1759), .B2(
        R2_SB_n361), .ZN(R2_SB_n396) );
  NAND2_X1 R2_SB_U370 ( .A1(R2_SB_n396), .A2(R2_SB_n397), .ZN(R2_SB_U8_Z_3) );
  AOI22_X1 R2_SB_U369 ( .A1(R2_n1726), .A2(R2_SB_n363), .B1(R2_n1694), .B2(
        R2_SB_n616), .ZN(R2_SB_n399) );
  AOI22_X1 R2_SB_U368 ( .A1(R2_n1662), .A2(R2_SB_n615), .B1(R2_n1758), .B2(
        R2_SB_n361), .ZN(R2_SB_n398) );
  NAND2_X1 R2_SB_U367 ( .A1(R2_SB_n398), .A2(R2_SB_n399), .ZN(R2_SB_U8_Z_2) );
  AOI22_X1 R2_SB_U366 ( .A1(R2_n1725), .A2(R2_SB_n363), .B1(R2_n1693), .B2(
        R2_SB_n616), .ZN(R2_SB_n401) );
  AOI22_X1 R2_SB_U365 ( .A1(R2_n1661), .A2(R2_SB_n615), .B1(R2_n1757), .B2(
        R2_SB_n361), .ZN(R2_SB_n400) );
  NAND2_X1 R2_SB_U364 ( .A1(R2_SB_n400), .A2(R2_SB_n401), .ZN(R2_SB_U8_Z_1) );
  AOI22_X1 R2_SB_U363 ( .A1(R2_n1724), .A2(R2_SB_n363), .B1(R2_n1692), .B2(
        R2_SB_n616), .ZN(R2_SB_n403) );
  AOI22_X1 R2_SB_U362 ( .A1(R2_n1660), .A2(R2_SB_n615), .B1(R2_n1756), .B2(
        R2_SB_n361), .ZN(R2_SB_n402) );
  NAND2_X1 R2_SB_U361 ( .A1(R2_SB_n402), .A2(R2_SB_n403), .ZN(R2_SB_U8_Z_0) );
  AOI22_X1 R2_SB_U360 ( .A1(R2_n1723), .A2(R2_SB_n363), .B1(R2_n1691), .B2(
        R2_SB_n616), .ZN(R2_SB_n372) );
  AOI22_X1 R2_SB_U359 ( .A1(R2_n1659), .A2(R2_SB_n615), .B1(R2_n1755), .B2(
        R2_SB_n361), .ZN(R2_SB_n371) );
  NAND2_X1 R2_SB_U358 ( .A1(R2_SB_n371), .A2(R2_SB_n372), .ZN(R2_SB_U9_Z_7) );
  AOI22_X1 R2_SB_U357 ( .A1(R2_n1722), .A2(R2_SB_n363), .B1(R2_n1690), .B2(
        R2_SB_n616), .ZN(R2_SB_n375) );
  AOI22_X1 R2_SB_U356 ( .A1(R2_n1658), .A2(R2_SB_n614), .B1(R2_n1754), .B2(
        R2_SB_n361), .ZN(R2_SB_n374) );
  NAND2_X1 R2_SB_U355 ( .A1(R2_SB_n374), .A2(R2_SB_n375), .ZN(R2_SB_U9_Z_6) );
  AOI22_X1 R2_SB_U354 ( .A1(R2_n1721), .A2(R2_SB_n363), .B1(R2_n1689), .B2(
        R2_SB_n616), .ZN(R2_SB_n377) );
  AOI22_X1 R2_SB_U353 ( .A1(R2_n1657), .A2(R2_SB_n614), .B1(R2_n1753), .B2(
        R2_SB_n361), .ZN(R2_SB_n376) );
  NAND2_X1 R2_SB_U352 ( .A1(R2_SB_n376), .A2(R2_SB_n377), .ZN(R2_SB_U9_Z_5) );
  AOI22_X1 R2_SB_U351 ( .A1(R2_n1720), .A2(R2_SB_n363), .B1(R2_n1688), .B2(
        R2_SB_n616), .ZN(R2_SB_n379) );
  AOI22_X1 R2_SB_U350 ( .A1(R2_n1656), .A2(R2_SB_n614), .B1(R2_n1752), .B2(
        R2_SB_n361), .ZN(R2_SB_n378) );
  NAND2_X1 R2_SB_U349 ( .A1(R2_SB_n378), .A2(R2_SB_n379), .ZN(R2_SB_U9_Z_4) );
  AOI22_X1 R2_SB_U348 ( .A1(R2_n1719), .A2(R2_SB_n363), .B1(R2_n1687), .B2(
        R2_SB_n616), .ZN(R2_SB_n381) );
  AOI22_X1 R2_SB_U347 ( .A1(R2_n1655), .A2(R2_SB_n614), .B1(R2_n1751), .B2(
        R2_SB_n361), .ZN(R2_SB_n380) );
  NAND2_X1 R2_SB_U346 ( .A1(R2_SB_n380), .A2(R2_SB_n381), .ZN(R2_SB_U9_Z_3) );
  AOI22_X1 R2_SB_U345 ( .A1(R2_n1718), .A2(R2_SB_n363), .B1(R2_n1686), .B2(
        R2_SB_n616), .ZN(R2_SB_n383) );
  AOI22_X1 R2_SB_U344 ( .A1(R2_n1654), .A2(R2_SB_n614), .B1(R2_n1750), .B2(
        R2_SB_n361), .ZN(R2_SB_n382) );
  NAND2_X1 R2_SB_U343 ( .A1(R2_SB_n382), .A2(R2_SB_n383), .ZN(R2_SB_U9_Z_2) );
  AOI22_X1 R2_SB_U342 ( .A1(R2_n1717), .A2(R2_SB_n617), .B1(R2_n1685), .B2(
        R2_SB_n616), .ZN(R2_SB_n385) );
  AOI22_X1 R2_SB_U341 ( .A1(R2_n1653), .A2(R2_SB_n614), .B1(R2_n1749), .B2(
        R2_SB_n361), .ZN(R2_SB_n384) );
  NAND2_X1 R2_SB_U340 ( .A1(R2_SB_n384), .A2(R2_SB_n385), .ZN(R2_SB_U9_Z_1) );
  AOI22_X1 R2_SB_U339 ( .A1(R2_n1716), .A2(R2_SB_n363), .B1(R2_n1684), .B2(
        R2_SB_n616), .ZN(R2_SB_n387) );
  AOI22_X1 R2_SB_U338 ( .A1(R2_n1652), .A2(R2_SB_n614), .B1(R2_n1748), .B2(
        R2_SB_n361), .ZN(R2_SB_n386) );
  NAND2_X1 R2_SB_U337 ( .A1(R2_SB_n386), .A2(R2_SB_n387), .ZN(R2_SB_U9_Z_0) );
  AOI22_X1 R2_SB_U336 ( .A1(R2_n1708), .A2(R2_SB_n617), .B1(R2_n1676), .B2(
        R2_SB_n367), .ZN(R2_SB_n441) );
  AOI22_X1 R2_SB_U335 ( .A1(R2_n1644), .A2(R2_SB_n614), .B1(R2_n1740), .B2(
        R2_SB_n618), .ZN(R2_SB_n440) );
  NAND2_X1 R2_SB_U334 ( .A1(R2_SB_n440), .A2(R2_SB_n441), .ZN(R2_SB_U10_Z_0)
         );
  XNOR2_X1 R2_SB_U333 ( .A(R2_SB_add_108_A_1_), .B(R2_SB_add_108_A_0_), .ZN(
        R2_SB_n425) );
  NOR2_X1 R2_SB_U332 ( .A1(R2_n1514), .A2(R2_SB_n425), .ZN(R2_SB_U4_Z_1) );
  OAI21_X1 R2_SB_U331 ( .B1(R2_SB_add_108_A_2_), .B2(R2_n1514), .A(R2_SB_n424), 
        .ZN(R2_SB_n421) );
  NOR3_X1 R2_SB_U330 ( .A1(R2_SB_n423), .A2(R2_SB_add_108_A_3_), .A3(R2_SB_n35), .ZN(R2_SB_n422) );
  AOI21_X1 R2_SB_U329 ( .B1(R2_SB_n421), .B2(R2_SB_add_108_A_3_), .A(
        R2_SB_n422), .ZN(R2_SB_n420) );
  INV_X1 R2_SB_U328 ( .A(R2_SB_n420), .ZN(R2_SB_n33) );
  NAND2_X1 R2_SB_U327 ( .A1(R2_SB_n144), .A2(R2_SB_n623), .ZN(R2_SB_n42) );
  OAI21_X1 R2_SB_U326 ( .B1(R2_SB_n32), .B2(R2_SB_n624), .A(R2_SB_n42), .ZN(
        R2_SB_n444) );
  NAND2_X1 R2_SB_U325 ( .A1(R2_SB_n80), .A2(R2_SB_n621), .ZN(R2_SB_n44) );
  OAI21_X1 R2_SB_U324 ( .B1(R2_SB_n32), .B2(R2_SB_n43), .A(R2_SB_n44), .ZN(
        R2_SB_n445) );
  NAND2_X1 R2_SB_U323 ( .A1(R2_SB_n112), .A2(R2_SB_n619), .ZN(R2_SB_n46) );
  OAI21_X1 R2_SB_U322 ( .B1(R2_SB_n32), .B2(R2_SB_n619), .A(R2_SB_n46), .ZN(
        R2_SB_n446) );
  NAND2_X1 R2_SB_U321 ( .A1(R2_SB_n176), .A2(R2_SB_n625), .ZN(R2_SB_n40) );
  OAI21_X1 R2_SB_U320 ( .B1(R2_SB_n39), .B2(R2_SB_n32), .A(R2_SB_n40), .ZN(
        R2_SB_n443) );
  NAND2_X1 R2_SB_U319 ( .A1(R2_SB_n169), .A2(R2_SB_n626), .ZN(R2_SB_n199) );
  OAI21_X1 R2_SB_U318 ( .B1(R2_SB_n39), .B2(R2_SB_n25), .A(R2_SB_n199), .ZN(
        R2_SB_n471) );
  NAND2_X1 R2_SB_U317 ( .A1(R2_SB_n137), .A2(R2_SB_n623), .ZN(R2_SB_n200) );
  OAI21_X1 R2_SB_U316 ( .B1(R2_SB_n624), .B2(R2_SB_n25), .A(R2_SB_n200), .ZN(
        R2_SB_n472) );
  NAND2_X1 R2_SB_U315 ( .A1(R2_SB_n73), .A2(R2_SB_n43), .ZN(R2_SB_n201) );
  OAI21_X1 R2_SB_U314 ( .B1(R2_SB_n621), .B2(R2_SB_n25), .A(R2_SB_n201), .ZN(
        R2_SB_n473) );
  NAND2_X1 R2_SB_U313 ( .A1(R2_SB_n105), .A2(R2_SB_n620), .ZN(R2_SB_n202) );
  OAI21_X1 R2_SB_U312 ( .B1(R2_SB_n45), .B2(R2_SB_n25), .A(R2_SB_n202), .ZN(
        R2_SB_n474) );
  NAND2_X1 R2_SB_U311 ( .A1(R2_SB_n173), .A2(R2_SB_n625), .ZN(R2_SB_n183) );
  OAI21_X1 R2_SB_U310 ( .B1(R2_SB_n626), .B2(R2_SB_n29), .A(R2_SB_n183), .ZN(
        R2_SB_n455) );
  NAND2_X1 R2_SB_U309 ( .A1(R2_SB_n141), .A2(R2_SB_n41), .ZN(R2_SB_n184) );
  OAI21_X1 R2_SB_U308 ( .B1(R2_SB_n623), .B2(R2_SB_n29), .A(R2_SB_n184), .ZN(
        R2_SB_n456) );
  NAND2_X1 R2_SB_U307 ( .A1(R2_SB_n77), .A2(R2_SB_n622), .ZN(R2_SB_n185) );
  OAI21_X1 R2_SB_U306 ( .B1(R2_SB_n43), .B2(R2_SB_n29), .A(R2_SB_n185), .ZN(
        R2_SB_n457) );
  NAND2_X1 R2_SB_U305 ( .A1(R2_SB_n109), .A2(R2_SB_n619), .ZN(R2_SB_n186) );
  OAI21_X1 R2_SB_U304 ( .B1(R2_SB_n620), .B2(R2_SB_n29), .A(R2_SB_n186), .ZN(
        R2_SB_n458) );
  NAND2_X1 R2_SB_U303 ( .A1(R2_SB_n174), .A2(R2_SB_n625), .ZN(R2_SB_n179) );
  OAI21_X1 R2_SB_U302 ( .B1(R2_SB_n39), .B2(R2_SB_n30), .A(R2_SB_n179), .ZN(
        R2_SB_n451) );
  NAND2_X1 R2_SB_U301 ( .A1(R2_SB_n142), .A2(R2_SB_n623), .ZN(R2_SB_n180) );
  OAI21_X1 R2_SB_U300 ( .B1(R2_SB_n624), .B2(R2_SB_n30), .A(R2_SB_n180), .ZN(
        R2_SB_n452) );
  NAND2_X1 R2_SB_U299 ( .A1(R2_SB_n78), .A2(R2_SB_n43), .ZN(R2_SB_n181) );
  OAI21_X1 R2_SB_U298 ( .B1(R2_SB_n622), .B2(R2_SB_n30), .A(R2_SB_n181), .ZN(
        R2_SB_n453) );
  NAND2_X1 R2_SB_U297 ( .A1(R2_SB_n110), .A2(R2_SB_n619), .ZN(R2_SB_n182) );
  OAI21_X1 R2_SB_U296 ( .B1(R2_SB_n45), .B2(R2_SB_n30), .A(R2_SB_n182), .ZN(
        R2_SB_n454) );
  NAND2_X1 R2_SB_U295 ( .A1(R2_SB_n175), .A2(R2_SB_n625), .ZN(R2_SB_n47) );
  OAI21_X1 R2_SB_U294 ( .B1(R2_SB_n626), .B2(R2_SB_n31), .A(R2_SB_n47), .ZN(
        R2_SB_n447) );
  NAND2_X1 R2_SB_U293 ( .A1(R2_SB_n143), .A2(R2_SB_n623), .ZN(R2_SB_n48) );
  OAI21_X1 R2_SB_U292 ( .B1(R2_SB_n623), .B2(R2_SB_n31), .A(R2_SB_n48), .ZN(
        R2_SB_n448) );
  NAND2_X1 R2_SB_U291 ( .A1(R2_SB_n79), .A2(R2_SB_n622), .ZN(R2_SB_n177) );
  OAI21_X1 R2_SB_U290 ( .B1(R2_SB_n43), .B2(R2_SB_n31), .A(R2_SB_n177), .ZN(
        R2_SB_n449) );
  NAND2_X1 R2_SB_U289 ( .A1(R2_SB_n111), .A2(R2_SB_n619), .ZN(R2_SB_n178) );
  OAI21_X1 R2_SB_U288 ( .B1(R2_SB_n620), .B2(R2_SB_n31), .A(R2_SB_n178), .ZN(
        R2_SB_n450) );
  NAND2_X1 R2_SB_U287 ( .A1(R2_SB_n161), .A2(R2_SB_n626), .ZN(R2_SB_n231) );
  OAI21_X1 R2_SB_U286 ( .B1(R2_SB_n39), .B2(R2_SB_n17), .A(R2_SB_n231), .ZN(
        R2_SB_n503) );
  NAND2_X1 R2_SB_U285 ( .A1(R2_SB_n129), .A2(R2_SB_n623), .ZN(R2_SB_n232) );
  OAI21_X1 R2_SB_U284 ( .B1(R2_SB_n41), .B2(R2_SB_n17), .A(R2_SB_n232), .ZN(
        R2_SB_n504) );
  NAND2_X1 R2_SB_U283 ( .A1(R2_SB_n65), .A2(R2_SB_n43), .ZN(R2_SB_n233) );
  OAI21_X1 R2_SB_U282 ( .B1(R2_SB_n621), .B2(R2_SB_n17), .A(R2_SB_n233), .ZN(
        R2_SB_n505) );
  NAND2_X1 R2_SB_U281 ( .A1(R2_SB_n97), .A2(R2_SB_n620), .ZN(R2_SB_n234) );
  OAI21_X1 R2_SB_U280 ( .B1(R2_SB_n45), .B2(R2_SB_n17), .A(R2_SB_n234), .ZN(
        R2_SB_n506) );
  NAND2_X1 R2_SB_U279 ( .A1(R2_SB_n163), .A2(R2_SB_n39), .ZN(R2_SB_n223) );
  OAI21_X1 R2_SB_U278 ( .B1(R2_SB_n39), .B2(R2_SB_n19), .A(R2_SB_n223), .ZN(
        R2_SB_n495) );
  NAND2_X1 R2_SB_U277 ( .A1(R2_SB_n131), .A2(R2_SB_n623), .ZN(R2_SB_n224) );
  OAI21_X1 R2_SB_U276 ( .B1(R2_SB_n624), .B2(R2_SB_n19), .A(R2_SB_n224), .ZN(
        R2_SB_n496) );
  NAND2_X1 R2_SB_U275 ( .A1(R2_SB_n67), .A2(R2_SB_n622), .ZN(R2_SB_n225) );
  OAI21_X1 R2_SB_U274 ( .B1(R2_SB_n621), .B2(R2_SB_n19), .A(R2_SB_n225), .ZN(
        R2_SB_n497) );
  NAND2_X1 R2_SB_U273 ( .A1(R2_SB_n99), .A2(R2_SB_n620), .ZN(R2_SB_n226) );
  OAI21_X1 R2_SB_U272 ( .B1(R2_SB_n45), .B2(R2_SB_n19), .A(R2_SB_n226), .ZN(
        R2_SB_n498) );
  NAND2_X1 R2_SB_U271 ( .A1(R2_SB_n165), .A2(R2_SB_n626), .ZN(R2_SB_n215) );
  OAI21_X1 R2_SB_U270 ( .B1(R2_SB_n626), .B2(R2_SB_n21), .A(R2_SB_n215), .ZN(
        R2_SB_n487) );
  NAND2_X1 R2_SB_U269 ( .A1(R2_SB_n133), .A2(R2_SB_n623), .ZN(R2_SB_n216) );
  OAI21_X1 R2_SB_U268 ( .B1(R2_SB_n624), .B2(R2_SB_n21), .A(R2_SB_n216), .ZN(
        R2_SB_n488) );
  NAND2_X1 R2_SB_U267 ( .A1(R2_SB_n69), .A2(R2_SB_n622), .ZN(R2_SB_n217) );
  OAI21_X1 R2_SB_U266 ( .B1(R2_SB_n622), .B2(R2_SB_n21), .A(R2_SB_n217), .ZN(
        R2_SB_n489) );
  NAND2_X1 R2_SB_U265 ( .A1(R2_SB_n101), .A2(R2_SB_n620), .ZN(R2_SB_n218) );
  OAI21_X1 R2_SB_U264 ( .B1(R2_SB_n45), .B2(R2_SB_n21), .A(R2_SB_n218), .ZN(
        R2_SB_n490) );
  NAND2_X1 R2_SB_U263 ( .A1(R2_SB_n168), .A2(R2_SB_n626), .ZN(R2_SB_n203) );
  OAI21_X1 R2_SB_U262 ( .B1(R2_SB_n625), .B2(R2_SB_n24), .A(R2_SB_n203), .ZN(
        R2_SB_n475) );
  NAND2_X1 R2_SB_U261 ( .A1(R2_SB_n134), .A2(R2_SB_n623), .ZN(R2_SB_n212) );
  OAI21_X1 R2_SB_U260 ( .B1(R2_SB_n624), .B2(R2_SB_n22), .A(R2_SB_n212), .ZN(
        R2_SB_n484) );
  NAND2_X1 R2_SB_U259 ( .A1(R2_SB_n70), .A2(R2_SB_n622), .ZN(R2_SB_n213) );
  OAI21_X1 R2_SB_U258 ( .B1(R2_SB_n43), .B2(R2_SB_n22), .A(R2_SB_n213), .ZN(
        R2_SB_n485) );
  NAND2_X1 R2_SB_U257 ( .A1(R2_SB_n102), .A2(R2_SB_n620), .ZN(R2_SB_n214) );
  OAI21_X1 R2_SB_U256 ( .B1(R2_SB_n45), .B2(R2_SB_n22), .A(R2_SB_n214), .ZN(
        R2_SB_n486) );
  NAND2_X1 R2_SB_U255 ( .A1(R2_SB_n167), .A2(R2_SB_n626), .ZN(R2_SB_n207) );
  OAI21_X1 R2_SB_U254 ( .B1(R2_SB_n626), .B2(R2_SB_n23), .A(R2_SB_n207), .ZN(
        R2_SB_n479) );
  NAND2_X1 R2_SB_U253 ( .A1(R2_SB_n135), .A2(R2_SB_n623), .ZN(R2_SB_n208) );
  OAI21_X1 R2_SB_U252 ( .B1(R2_SB_n624), .B2(R2_SB_n23), .A(R2_SB_n208), .ZN(
        R2_SB_n480) );
  NAND2_X1 R2_SB_U251 ( .A1(R2_SB_n71), .A2(R2_SB_n622), .ZN(R2_SB_n209) );
  OAI21_X1 R2_SB_U250 ( .B1(R2_SB_n43), .B2(R2_SB_n23), .A(R2_SB_n209), .ZN(
        R2_SB_n481) );
  NAND2_X1 R2_SB_U249 ( .A1(R2_SB_n103), .A2(R2_SB_n620), .ZN(R2_SB_n210) );
  OAI21_X1 R2_SB_U248 ( .B1(R2_SB_n45), .B2(R2_SB_n23), .A(R2_SB_n210), .ZN(
        R2_SB_n482) );
  NAND2_X1 R2_SB_U247 ( .A1(R2_SB_n136), .A2(R2_SB_n623), .ZN(R2_SB_n204) );
  OAI21_X1 R2_SB_U246 ( .B1(R2_SB_n624), .B2(R2_SB_n24), .A(R2_SB_n204), .ZN(
        R2_SB_n476) );
  NAND2_X1 R2_SB_U245 ( .A1(R2_SB_n72), .A2(R2_SB_n622), .ZN(R2_SB_n205) );
  OAI21_X1 R2_SB_U244 ( .B1(R2_SB_n43), .B2(R2_SB_n24), .A(R2_SB_n205), .ZN(
        R2_SB_n477) );
  NAND2_X1 R2_SB_U243 ( .A1(R2_SB_n104), .A2(R2_SB_n620), .ZN(R2_SB_n206) );
  OAI21_X1 R2_SB_U242 ( .B1(R2_SB_n45), .B2(R2_SB_n24), .A(R2_SB_n206), .ZN(
        R2_SB_n478) );
  NAND2_X1 R2_SB_U241 ( .A1(R2_SB_n153), .A2(R2_SB_n39), .ZN(R2_SB_n263) );
  OAI21_X1 R2_SB_U240 ( .B1(R2_SB_n39), .B2(R2_SB_n9), .A(R2_SB_n263), .ZN(
        R2_SB_n535) );
  NAND2_X1 R2_SB_U239 ( .A1(R2_SB_n121), .A2(R2_SB_n41), .ZN(R2_SB_n264) );
  OAI21_X1 R2_SB_U238 ( .B1(R2_SB_n41), .B2(R2_SB_n9), .A(R2_SB_n264), .ZN(
        R2_SB_n536) );
  NAND2_X1 R2_SB_U237 ( .A1(R2_SB_n57), .A2(R2_SB_n622), .ZN(R2_SB_n265) );
  OAI21_X1 R2_SB_U236 ( .B1(R2_SB_n621), .B2(R2_SB_n9), .A(R2_SB_n265), .ZN(
        R2_SB_n537) );
  NAND2_X1 R2_SB_U235 ( .A1(R2_SB_n89), .A2(R2_SB_n619), .ZN(R2_SB_n266) );
  OAI21_X1 R2_SB_U234 ( .B1(R2_SB_n619), .B2(R2_SB_n9), .A(R2_SB_n266), .ZN(
        R2_SB_n538) );
  NAND2_X1 R2_SB_U233 ( .A1(R2_SB_n155), .A2(R2_SB_n39), .ZN(R2_SB_n255) );
  OAI21_X1 R2_SB_U232 ( .B1(R2_SB_n39), .B2(R2_SB_n11), .A(R2_SB_n255), .ZN(
        R2_SB_n527) );
  NAND2_X1 R2_SB_U231 ( .A1(R2_SB_n123), .A2(R2_SB_n41), .ZN(R2_SB_n256) );
  OAI21_X1 R2_SB_U230 ( .B1(R2_SB_n41), .B2(R2_SB_n11), .A(R2_SB_n256), .ZN(
        R2_SB_n528) );
  NAND2_X1 R2_SB_U229 ( .A1(R2_SB_n59), .A2(R2_SB_n622), .ZN(R2_SB_n257) );
  OAI21_X1 R2_SB_U228 ( .B1(R2_SB_n621), .B2(R2_SB_n11), .A(R2_SB_n257), .ZN(
        R2_SB_n529) );
  NAND2_X1 R2_SB_U227 ( .A1(R2_SB_n91), .A2(R2_SB_n619), .ZN(R2_SB_n258) );
  OAI21_X1 R2_SB_U226 ( .B1(R2_SB_n620), .B2(R2_SB_n11), .A(R2_SB_n258), .ZN(
        R2_SB_n530) );
  NAND2_X1 R2_SB_U225 ( .A1(R2_SB_n157), .A2(R2_SB_n39), .ZN(R2_SB_n247) );
  OAI21_X1 R2_SB_U224 ( .B1(R2_SB_n39), .B2(R2_SB_n13), .A(R2_SB_n247), .ZN(
        R2_SB_n519) );
  NAND2_X1 R2_SB_U223 ( .A1(R2_SB_n125), .A2(R2_SB_n41), .ZN(R2_SB_n248) );
  OAI21_X1 R2_SB_U222 ( .B1(R2_SB_n41), .B2(R2_SB_n13), .A(R2_SB_n248), .ZN(
        R2_SB_n520) );
  NAND2_X1 R2_SB_U221 ( .A1(R2_SB_n61), .A2(R2_SB_n622), .ZN(R2_SB_n249) );
  OAI21_X1 R2_SB_U220 ( .B1(R2_SB_n621), .B2(R2_SB_n13), .A(R2_SB_n249), .ZN(
        R2_SB_n521) );
  NAND2_X1 R2_SB_U219 ( .A1(R2_SB_n93), .A2(R2_SB_n45), .ZN(R2_SB_n250) );
  OAI21_X1 R2_SB_U218 ( .B1(R2_SB_n45), .B2(R2_SB_n13), .A(R2_SB_n250), .ZN(
        R2_SB_n522) );
  NAND2_X1 R2_SB_U217 ( .A1(R2_SB_n158), .A2(R2_SB_n39), .ZN(R2_SB_n243) );
  OAI21_X1 R2_SB_U216 ( .B1(R2_SB_n39), .B2(R2_SB_n14), .A(R2_SB_n243), .ZN(
        R2_SB_n515) );
  NAND2_X1 R2_SB_U215 ( .A1(R2_SB_n126), .A2(R2_SB_n41), .ZN(R2_SB_n244) );
  OAI21_X1 R2_SB_U214 ( .B1(R2_SB_n41), .B2(R2_SB_n14), .A(R2_SB_n244), .ZN(
        R2_SB_n516) );
  NAND2_X1 R2_SB_U213 ( .A1(R2_SB_n62), .A2(R2_SB_n622), .ZN(R2_SB_n245) );
  OAI21_X1 R2_SB_U212 ( .B1(R2_SB_n621), .B2(R2_SB_n14), .A(R2_SB_n245), .ZN(
        R2_SB_n517) );
  NAND2_X1 R2_SB_U211 ( .A1(R2_SB_n94), .A2(R2_SB_n45), .ZN(R2_SB_n246) );
  OAI21_X1 R2_SB_U210 ( .B1(R2_SB_n45), .B2(R2_SB_n14), .A(R2_SB_n246), .ZN(
        R2_SB_n518) );
  NAND2_X1 R2_SB_U209 ( .A1(R2_SB_n159), .A2(R2_SB_n39), .ZN(R2_SB_n239) );
  OAI21_X1 R2_SB_U208 ( .B1(R2_SB_n39), .B2(R2_SB_n15), .A(R2_SB_n239), .ZN(
        R2_SB_n511) );
  NAND2_X1 R2_SB_U207 ( .A1(R2_SB_n127), .A2(R2_SB_n41), .ZN(R2_SB_n240) );
  OAI21_X1 R2_SB_U206 ( .B1(R2_SB_n41), .B2(R2_SB_n15), .A(R2_SB_n240), .ZN(
        R2_SB_n512) );
  NAND2_X1 R2_SB_U205 ( .A1(R2_SB_n63), .A2(R2_SB_n622), .ZN(R2_SB_n241) );
  OAI21_X1 R2_SB_U204 ( .B1(R2_SB_n621), .B2(R2_SB_n15), .A(R2_SB_n241), .ZN(
        R2_SB_n513) );
  NAND2_X1 R2_SB_U203 ( .A1(R2_SB_n95), .A2(R2_SB_n45), .ZN(R2_SB_n242) );
  OAI21_X1 R2_SB_U202 ( .B1(R2_SB_n45), .B2(R2_SB_n15), .A(R2_SB_n242), .ZN(
        R2_SB_n514) );
  NAND2_X1 R2_SB_U201 ( .A1(R2_SB_n160), .A2(R2_SB_n625), .ZN(R2_SB_n235) );
  OAI21_X1 R2_SB_U200 ( .B1(R2_SB_n39), .B2(R2_SB_n16), .A(R2_SB_n235), .ZN(
        R2_SB_n507) );
  NAND2_X1 R2_SB_U199 ( .A1(R2_SB_n128), .A2(R2_SB_n41), .ZN(R2_SB_n236) );
  OAI21_X1 R2_SB_U198 ( .B1(R2_SB_n41), .B2(R2_SB_n16), .A(R2_SB_n236), .ZN(
        R2_SB_n508) );
  NAND2_X1 R2_SB_U197 ( .A1(R2_SB_n64), .A2(R2_SB_n622), .ZN(R2_SB_n237) );
  OAI21_X1 R2_SB_U196 ( .B1(R2_SB_n621), .B2(R2_SB_n16), .A(R2_SB_n237), .ZN(
        R2_SB_n509) );
  NAND2_X1 R2_SB_U195 ( .A1(R2_SB_n96), .A2(R2_SB_n45), .ZN(R2_SB_n238) );
  OAI21_X1 R2_SB_U194 ( .B1(R2_SB_n45), .B2(R2_SB_n16), .A(R2_SB_n238), .ZN(
        R2_SB_n510) );
  NAND2_X1 R2_SB_U193 ( .A1(R2_SB_n145), .A2(R2_SB_n625), .ZN(R2_SB_n360) );
  OAI21_X1 R2_SB_U192 ( .B1(R2_SB_n626), .B2(R2_SB_n1), .A(R2_SB_n360), .ZN(
        R2_SB_n567) );
  NAND2_X1 R2_SB_U191 ( .A1(R2_SB_n113), .A2(R2_SB_n623), .ZN(R2_SB_n362) );
  OAI21_X1 R2_SB_U190 ( .B1(R2_SB_n623), .B2(R2_SB_n1), .A(R2_SB_n362), .ZN(
        R2_SB_n568) );
  NAND2_X1 R2_SB_U189 ( .A1(R2_SB_n49), .A2(R2_SB_n43), .ZN(R2_SB_n364) );
  OAI21_X1 R2_SB_U188 ( .B1(R2_SB_n43), .B2(R2_SB_n1), .A(R2_SB_n364), .ZN(
        R2_SB_n569) );
  NAND2_X1 R2_SB_U187 ( .A1(R2_SB_n81), .A2(R2_SB_n619), .ZN(R2_SB_n366) );
  OAI21_X1 R2_SB_U186 ( .B1(R2_SB_n620), .B2(R2_SB_n1), .A(R2_SB_n366), .ZN(
        R2_SB_n570) );
  NAND2_X1 R2_SB_U185 ( .A1(R2_SB_n147), .A2(R2_SB_n625), .ZN(R2_SB_n352) );
  OAI21_X1 R2_SB_U184 ( .B1(R2_SB_n625), .B2(R2_SB_n3), .A(R2_SB_n352), .ZN(
        R2_SB_n559) );
  NAND2_X1 R2_SB_U183 ( .A1(R2_SB_n115), .A2(R2_SB_n623), .ZN(R2_SB_n353) );
  OAI21_X1 R2_SB_U182 ( .B1(R2_SB_n624), .B2(R2_SB_n3), .A(R2_SB_n353), .ZN(
        R2_SB_n560) );
  NAND2_X1 R2_SB_U181 ( .A1(R2_SB_n51), .A2(R2_SB_n43), .ZN(R2_SB_n354) );
  OAI21_X1 R2_SB_U180 ( .B1(R2_SB_n43), .B2(R2_SB_n3), .A(R2_SB_n354), .ZN(
        R2_SB_n561) );
  NAND2_X1 R2_SB_U179 ( .A1(R2_SB_n83), .A2(R2_SB_n619), .ZN(R2_SB_n355) );
  OAI21_X1 R2_SB_U178 ( .B1(R2_SB_n45), .B2(R2_SB_n3), .A(R2_SB_n355), .ZN(
        R2_SB_n562) );
  NAND2_X1 R2_SB_U177 ( .A1(R2_SB_n149), .A2(R2_SB_n625), .ZN(R2_SB_n280) );
  OAI21_X1 R2_SB_U176 ( .B1(R2_SB_n39), .B2(R2_SB_n5), .A(R2_SB_n280), .ZN(
        R2_SB_n551) );
  NAND2_X1 R2_SB_U175 ( .A1(R2_SB_n117), .A2(R2_SB_n623), .ZN(R2_SB_n345) );
  OAI21_X1 R2_SB_U174 ( .B1(R2_SB_n41), .B2(R2_SB_n5), .A(R2_SB_n345), .ZN(
        R2_SB_n552) );
  NAND2_X1 R2_SB_U173 ( .A1(R2_SB_n53), .A2(R2_SB_n43), .ZN(R2_SB_n346) );
  OAI21_X1 R2_SB_U172 ( .B1(R2_SB_n621), .B2(R2_SB_n5), .A(R2_SB_n346), .ZN(
        R2_SB_n553) );
  NAND2_X1 R2_SB_U171 ( .A1(R2_SB_n85), .A2(R2_SB_n619), .ZN(R2_SB_n347) );
  OAI21_X1 R2_SB_U170 ( .B1(R2_SB_n45), .B2(R2_SB_n5), .A(R2_SB_n347), .ZN(
        R2_SB_n554) );
  NAND2_X1 R2_SB_U169 ( .A1(R2_SB_n150), .A2(R2_SB_n625), .ZN(R2_SB_n275) );
  OAI21_X1 R2_SB_U168 ( .B1(R2_SB_n39), .B2(R2_SB_n6), .A(R2_SB_n275), .ZN(
        R2_SB_n547) );
  NAND2_X1 R2_SB_U167 ( .A1(R2_SB_n118), .A2(R2_SB_n41), .ZN(R2_SB_n277) );
  OAI21_X1 R2_SB_U166 ( .B1(R2_SB_n41), .B2(R2_SB_n6), .A(R2_SB_n277), .ZN(
        R2_SB_n548) );
  NAND2_X1 R2_SB_U165 ( .A1(R2_SB_n54), .A2(R2_SB_n621), .ZN(R2_SB_n278) );
  OAI21_X1 R2_SB_U164 ( .B1(R2_SB_n621), .B2(R2_SB_n6), .A(R2_SB_n278), .ZN(
        R2_SB_n549) );
  NAND2_X1 R2_SB_U163 ( .A1(R2_SB_n86), .A2(R2_SB_n620), .ZN(R2_SB_n279) );
  OAI21_X1 R2_SB_U162 ( .B1(R2_SB_n45), .B2(R2_SB_n6), .A(R2_SB_n279), .ZN(
        R2_SB_n550) );
  NAND2_X1 R2_SB_U161 ( .A1(R2_SB_n151), .A2(R2_SB_n625), .ZN(R2_SB_n271) );
  OAI21_X1 R2_SB_U160 ( .B1(R2_SB_n39), .B2(R2_SB_n7), .A(R2_SB_n271), .ZN(
        R2_SB_n543) );
  NAND2_X1 R2_SB_U159 ( .A1(R2_SB_n119), .A2(R2_SB_n41), .ZN(R2_SB_n272) );
  OAI21_X1 R2_SB_U158 ( .B1(R2_SB_n41), .B2(R2_SB_n7), .A(R2_SB_n272), .ZN(
        R2_SB_n544) );
  NAND2_X1 R2_SB_U157 ( .A1(R2_SB_n55), .A2(R2_SB_n43), .ZN(R2_SB_n273) );
  OAI21_X1 R2_SB_U156 ( .B1(R2_SB_n621), .B2(R2_SB_n7), .A(R2_SB_n273), .ZN(
        R2_SB_n545) );
  NAND2_X1 R2_SB_U155 ( .A1(R2_SB_n87), .A2(R2_SB_n619), .ZN(R2_SB_n274) );
  OAI21_X1 R2_SB_U154 ( .B1(R2_SB_n619), .B2(R2_SB_n7), .A(R2_SB_n274), .ZN(
        R2_SB_n546) );
  NAND2_X1 R2_SB_U153 ( .A1(R2_SB_n152), .A2(R2_SB_n625), .ZN(R2_SB_n267) );
  OAI21_X1 R2_SB_U152 ( .B1(R2_SB_n626), .B2(R2_SB_n8), .A(R2_SB_n267), .ZN(
        R2_SB_n539) );
  NAND2_X1 R2_SB_U151 ( .A1(R2_SB_n120), .A2(R2_SB_n623), .ZN(R2_SB_n268) );
  OAI21_X1 R2_SB_U150 ( .B1(R2_SB_n41), .B2(R2_SB_n8), .A(R2_SB_n268), .ZN(
        R2_SB_n540) );
  NAND2_X1 R2_SB_U149 ( .A1(R2_SB_n56), .A2(R2_SB_n621), .ZN(R2_SB_n269) );
  OAI21_X1 R2_SB_U148 ( .B1(R2_SB_n621), .B2(R2_SB_n8), .A(R2_SB_n269), .ZN(
        R2_SB_n541) );
  NAND2_X1 R2_SB_U147 ( .A1(R2_SB_n88), .A2(R2_SB_n619), .ZN(R2_SB_n270) );
  OAI21_X1 R2_SB_U146 ( .B1(R2_SB_n619), .B2(R2_SB_n8), .A(R2_SB_n270), .ZN(
        R2_SB_n542) );
  NAND2_X1 R2_SB_U145 ( .A1(R2_SB_n171), .A2(R2_SB_n626), .ZN(R2_SB_n191) );
  OAI21_X1 R2_SB_U144 ( .B1(R2_SB_n39), .B2(R2_SB_n27), .A(R2_SB_n191), .ZN(
        R2_SB_n463) );
  NAND2_X1 R2_SB_U143 ( .A1(R2_SB_n139), .A2(R2_SB_n41), .ZN(R2_SB_n192) );
  OAI21_X1 R2_SB_U142 ( .B1(R2_SB_n624), .B2(R2_SB_n27), .A(R2_SB_n192), .ZN(
        R2_SB_n464) );
  NAND2_X1 R2_SB_U141 ( .A1(R2_SB_n75), .A2(R2_SB_n622), .ZN(R2_SB_n193) );
  OAI21_X1 R2_SB_U140 ( .B1(R2_SB_n43), .B2(R2_SB_n27), .A(R2_SB_n193), .ZN(
        R2_SB_n465) );
  NAND2_X1 R2_SB_U139 ( .A1(R2_SB_n107), .A2(R2_SB_n45), .ZN(R2_SB_n194) );
  OAI21_X1 R2_SB_U138 ( .B1(R2_SB_n45), .B2(R2_SB_n27), .A(R2_SB_n194), .ZN(
        R2_SB_n466) );
  NAND2_X1 R2_SB_U137 ( .A1(R2_SB_n166), .A2(R2_SB_n626), .ZN(R2_SB_n211) );
  OAI21_X1 R2_SB_U136 ( .B1(R2_SB_n625), .B2(R2_SB_n22), .A(R2_SB_n211), .ZN(
        R2_SB_n483) );
  NAND2_X1 R2_SB_U135 ( .A1(R2_SB_n170), .A2(R2_SB_n626), .ZN(R2_SB_n195) );
  OAI21_X1 R2_SB_U134 ( .B1(R2_SB_n625), .B2(R2_SB_n26), .A(R2_SB_n195), .ZN(
        R2_SB_n467) );
  NAND2_X1 R2_SB_U133 ( .A1(R2_SB_n138), .A2(R2_SB_n41), .ZN(R2_SB_n196) );
  OAI21_X1 R2_SB_U132 ( .B1(R2_SB_n624), .B2(R2_SB_n26), .A(R2_SB_n196), .ZN(
        R2_SB_n468) );
  NAND2_X1 R2_SB_U131 ( .A1(R2_SB_n74), .A2(R2_SB_n622), .ZN(R2_SB_n197) );
  OAI21_X1 R2_SB_U130 ( .B1(R2_SB_n43), .B2(R2_SB_n26), .A(R2_SB_n197), .ZN(
        R2_SB_n469) );
  NAND2_X1 R2_SB_U129 ( .A1(R2_SB_n106), .A2(R2_SB_n619), .ZN(R2_SB_n198) );
  OAI21_X1 R2_SB_U128 ( .B1(R2_SB_n45), .B2(R2_SB_n26), .A(R2_SB_n198), .ZN(
        R2_SB_n470) );
  NAND2_X1 R2_SB_U127 ( .A1(R2_SB_n162), .A2(R2_SB_n626), .ZN(R2_SB_n227) );
  OAI21_X1 R2_SB_U126 ( .B1(R2_SB_n626), .B2(R2_SB_n18), .A(R2_SB_n227), .ZN(
        R2_SB_n499) );
  NAND2_X1 R2_SB_U125 ( .A1(R2_SB_n130), .A2(R2_SB_n623), .ZN(R2_SB_n228) );
  OAI21_X1 R2_SB_U124 ( .B1(R2_SB_n624), .B2(R2_SB_n18), .A(R2_SB_n228), .ZN(
        R2_SB_n500) );
  NAND2_X1 R2_SB_U123 ( .A1(R2_SB_n66), .A2(R2_SB_n622), .ZN(R2_SB_n229) );
  OAI21_X1 R2_SB_U122 ( .B1(R2_SB_n43), .B2(R2_SB_n18), .A(R2_SB_n229), .ZN(
        R2_SB_n501) );
  NAND2_X1 R2_SB_U121 ( .A1(R2_SB_n98), .A2(R2_SB_n620), .ZN(R2_SB_n230) );
  OAI21_X1 R2_SB_U120 ( .B1(R2_SB_n45), .B2(R2_SB_n18), .A(R2_SB_n230), .ZN(
        R2_SB_n502) );
  NAND2_X1 R2_SB_U119 ( .A1(R2_SB_n154), .A2(R2_SB_n39), .ZN(R2_SB_n259) );
  OAI21_X1 R2_SB_U118 ( .B1(R2_SB_n625), .B2(R2_SB_n10), .A(R2_SB_n259), .ZN(
        R2_SB_n531) );
  NAND2_X1 R2_SB_U117 ( .A1(R2_SB_n122), .A2(R2_SB_n41), .ZN(R2_SB_n260) );
  OAI21_X1 R2_SB_U116 ( .B1(R2_SB_n623), .B2(R2_SB_n10), .A(R2_SB_n260), .ZN(
        R2_SB_n532) );
  NAND2_X1 R2_SB_U115 ( .A1(R2_SB_n58), .A2(R2_SB_n622), .ZN(R2_SB_n261) );
  OAI21_X1 R2_SB_U114 ( .B1(R2_SB_n621), .B2(R2_SB_n10), .A(R2_SB_n261), .ZN(
        R2_SB_n533) );
  NAND2_X1 R2_SB_U113 ( .A1(R2_SB_n90), .A2(R2_SB_n619), .ZN(R2_SB_n262) );
  OAI21_X1 R2_SB_U112 ( .B1(R2_SB_n619), .B2(R2_SB_n10), .A(R2_SB_n262), .ZN(
        R2_SB_n534) );
  NAND2_X1 R2_SB_U111 ( .A1(R2_SB_n146), .A2(R2_SB_n625), .ZN(R2_SB_n356) );
  OAI21_X1 R2_SB_U110 ( .B1(R2_SB_n626), .B2(R2_SB_n2), .A(R2_SB_n356), .ZN(
        R2_SB_n563) );
  NAND2_X1 R2_SB_U109 ( .A1(R2_SB_n114), .A2(R2_SB_n623), .ZN(R2_SB_n357) );
  OAI21_X1 R2_SB_U108 ( .B1(R2_SB_n624), .B2(R2_SB_n2), .A(R2_SB_n357), .ZN(
        R2_SB_n564) );
  NAND2_X1 R2_SB_U107 ( .A1(R2_SB_n50), .A2(R2_SB_n43), .ZN(R2_SB_n358) );
  OAI21_X1 R2_SB_U106 ( .B1(R2_SB_n43), .B2(R2_SB_n2), .A(R2_SB_n358), .ZN(
        R2_SB_n565) );
  NAND2_X1 R2_SB_U105 ( .A1(R2_SB_n82), .A2(R2_SB_n619), .ZN(R2_SB_n359) );
  OAI21_X1 R2_SB_U104 ( .B1(R2_SB_n620), .B2(R2_SB_n2), .A(R2_SB_n359), .ZN(
        R2_SB_n566) );
  NAND2_X1 R2_SB_U103 ( .A1(R2_SB_n172), .A2(R2_SB_n626), .ZN(R2_SB_n187) );
  OAI21_X1 R2_SB_U102 ( .B1(R2_SB_n626), .B2(R2_SB_n28), .A(R2_SB_n187), .ZN(
        R2_SB_n459) );
  NAND2_X1 R2_SB_U101 ( .A1(R2_SB_n140), .A2(R2_SB_n623), .ZN(R2_SB_n188) );
  OAI21_X1 R2_SB_U100 ( .B1(R2_SB_n624), .B2(R2_SB_n28), .A(R2_SB_n188), .ZN(
        R2_SB_n460) );
  NAND2_X1 R2_SB_U99 ( .A1(R2_SB_n76), .A2(R2_SB_n622), .ZN(R2_SB_n189) );
  OAI21_X1 R2_SB_U98 ( .B1(R2_SB_n43), .B2(R2_SB_n28), .A(R2_SB_n189), .ZN(
        R2_SB_n461) );
  NAND2_X1 R2_SB_U97 ( .A1(R2_SB_n108), .A2(R2_SB_n620), .ZN(R2_SB_n190) );
  OAI21_X1 R2_SB_U96 ( .B1(R2_SB_n45), .B2(R2_SB_n28), .A(R2_SB_n190), .ZN(
        R2_SB_n462) );
  NAND2_X1 R2_SB_U95 ( .A1(R2_SB_n164), .A2(R2_SB_n626), .ZN(R2_SB_n219) );
  OAI21_X1 R2_SB_U94 ( .B1(R2_SB_n39), .B2(R2_SB_n20), .A(R2_SB_n219), .ZN(
        R2_SB_n491) );
  NAND2_X1 R2_SB_U93 ( .A1(R2_SB_n132), .A2(R2_SB_n623), .ZN(R2_SB_n220) );
  OAI21_X1 R2_SB_U92 ( .B1(R2_SB_n624), .B2(R2_SB_n20), .A(R2_SB_n220), .ZN(
        R2_SB_n492) );
  NAND2_X1 R2_SB_U91 ( .A1(R2_SB_n68), .A2(R2_SB_n622), .ZN(R2_SB_n221) );
  OAI21_X1 R2_SB_U90 ( .B1(R2_SB_n43), .B2(R2_SB_n20), .A(R2_SB_n221), .ZN(
        R2_SB_n493) );
  NAND2_X1 R2_SB_U89 ( .A1(R2_SB_n100), .A2(R2_SB_n620), .ZN(R2_SB_n222) );
  OAI21_X1 R2_SB_U88 ( .B1(R2_SB_n619), .B2(R2_SB_n20), .A(R2_SB_n222), .ZN(
        R2_SB_n494) );
  NAND2_X1 R2_SB_U87 ( .A1(R2_SB_n156), .A2(R2_SB_n625), .ZN(R2_SB_n251) );
  OAI21_X1 R2_SB_U86 ( .B1(R2_SB_n626), .B2(R2_SB_n12), .A(R2_SB_n251), .ZN(
        R2_SB_n523) );
  NAND2_X1 R2_SB_U85 ( .A1(R2_SB_n124), .A2(R2_SB_n41), .ZN(R2_SB_n252) );
  OAI21_X1 R2_SB_U84 ( .B1(R2_SB_n623), .B2(R2_SB_n12), .A(R2_SB_n252), .ZN(
        R2_SB_n524) );
  NAND2_X1 R2_SB_U83 ( .A1(R2_SB_n60), .A2(R2_SB_n622), .ZN(R2_SB_n253) );
  OAI21_X1 R2_SB_U82 ( .B1(R2_SB_n621), .B2(R2_SB_n12), .A(R2_SB_n253), .ZN(
        R2_SB_n525) );
  NAND2_X1 R2_SB_U81 ( .A1(R2_SB_n92), .A2(R2_SB_n619), .ZN(R2_SB_n254) );
  OAI21_X1 R2_SB_U80 ( .B1(R2_SB_n619), .B2(R2_SB_n12), .A(R2_SB_n254), .ZN(
        R2_SB_n526) );
  NAND2_X1 R2_SB_U79 ( .A1(R2_SB_n148), .A2(R2_SB_n625), .ZN(R2_SB_n348) );
  OAI21_X1 R2_SB_U78 ( .B1(R2_SB_n625), .B2(R2_SB_n4), .A(R2_SB_n348), .ZN(
        R2_SB_n555) );
  NAND2_X1 R2_SB_U77 ( .A1(R2_SB_n116), .A2(R2_SB_n623), .ZN(R2_SB_n349) );
  OAI21_X1 R2_SB_U76 ( .B1(R2_SB_n624), .B2(R2_SB_n4), .A(R2_SB_n349), .ZN(
        R2_SB_n556) );
  NAND2_X1 R2_SB_U75 ( .A1(R2_SB_n52), .A2(R2_SB_n621), .ZN(R2_SB_n350) );
  OAI21_X1 R2_SB_U74 ( .B1(R2_SB_n621), .B2(R2_SB_n4), .A(R2_SB_n350), .ZN(
        R2_SB_n557) );
  NAND2_X1 R2_SB_U73 ( .A1(R2_SB_n84), .A2(R2_SB_n619), .ZN(R2_SB_n351) );
  OAI21_X1 R2_SB_U72 ( .B1(R2_SB_n619), .B2(R2_SB_n4), .A(R2_SB_n351), .ZN(
        R2_SB_n558) );
  NAND2_X1 R2_SB_U71 ( .A1(R2_SB_n276), .A2(R2_SB_n368), .ZN(R2_SB_n369) );
  OAI21_X1 R2_SB_U70 ( .B1(R2_n1514), .B2(R2_SB_n368), .A(R2_SB_n369), .ZN(
        R2_SB_n571) );
  NAND2_X1 R2_SB_U69 ( .A1(R2_n1515), .A2(R2_SB_n368), .ZN(R2_SB_n370) );
  OAI21_X1 R2_SB_U68 ( .B1(R2_n1514), .B2(R2_SB_n368), .A(R2_SB_n370), .ZN(
        R2_SB_n572) );
  INV_X1 R2_SB_U67 ( .A(R2_n1514), .ZN(R2_SB_n38) );
  OAI22_X1 R2_SB_U66 ( .A1(R2_SB_n424), .A2(R2_SB_n35), .B1(R2_SB_add_108_A_2_), .B2(R2_SB_n423), .ZN(R2_SB_U4_Z_2) );
  NOR2_X1 R2_SB_U63 ( .A1(R2_SB_add_108_A_0_), .A2(R2_n1514), .ZN(R2_SB_U4_Z_0) );
  AOI21_X1 R2_SB_U62 ( .B1(R2_SB_n38), .B2(R2_SB_n36), .A(R2_SB_U4_Z_0), .ZN(
        R2_SB_n424) );
  NOR3_X1 R2_SB_U61 ( .A1(R2_SB_add_108_A_2_), .A2(R2_SB_add_108_A_3_), .A3(
        R2_SB_n36), .ZN(R2_SB_n442) );
  NOR3_X1 R2_SB_U59 ( .A1(R2_SB_add_108_A_2_), .A2(R2_SB_add_108_A_3_), .A3(
        R2_SB_add_108_A_1_), .ZN(R2_SB_n365) );
  NOR2_X1 R2_SB_U58 ( .A1(R2_n1514), .A2(R2_SB_n618), .ZN(R2_SB_n368) );
  INV_X1 R2_SB_U57 ( .A(R2_SB_n[288]), .ZN(R2_SB_n32) );
  INV_X1 R2_SB_U56 ( .A(R2_SB_n304), .ZN(R2_SB_n24) );
  INV_X1 R2_SB_U55 ( .A(R2_SB_n320), .ZN(R2_SB_n16) );
  INV_X1 R2_SB_U54 ( .A(R2_SB_n336), .ZN(R2_SB_n8) );
  INV_X1 R2_SB_U53 ( .A(R2_SB_n[281]), .ZN(R2_SB_n25) );
  INV_X1 R2_SB_U52 ( .A(R2_SB_n[283]), .ZN(R2_SB_n27) );
  INV_X1 R2_SB_U51 ( .A(R2_SB_n[284]), .ZN(R2_SB_n28) );
  INV_X1 R2_SB_U50 ( .A(R2_SB_n[285]), .ZN(R2_SB_n29) );
  INV_X1 R2_SB_U49 ( .A(R2_SB_n297), .ZN(R2_SB_n17) );
  INV_X1 R2_SB_U48 ( .A(R2_SB_n299), .ZN(R2_SB_n19) );
  INV_X1 R2_SB_U47 ( .A(R2_SB_n300), .ZN(R2_SB_n20) );
  INV_X1 R2_SB_U46 ( .A(R2_SB_n301), .ZN(R2_SB_n21) );
  INV_X1 R2_SB_U45 ( .A(R2_SB_n313), .ZN(R2_SB_n9) );
  INV_X1 R2_SB_U44 ( .A(R2_SB_n315), .ZN(R2_SB_n11) );
  INV_X1 R2_SB_U43 ( .A(R2_SB_n316), .ZN(R2_SB_n12) );
  INV_X1 R2_SB_U42 ( .A(R2_SB_n317), .ZN(R2_SB_n13) );
  INV_X1 R2_SB_U41 ( .A(R2_SB_n329), .ZN(R2_SB_n1) );
  INV_X1 R2_SB_U40 ( .A(R2_SB_n331), .ZN(R2_SB_n3) );
  INV_X1 R2_SB_U39 ( .A(R2_SB_n332), .ZN(R2_SB_n4) );
  INV_X1 R2_SB_U38 ( .A(R2_SB_n333), .ZN(R2_SB_n5) );
  INV_X1 R2_SB_U37 ( .A(R2_SB_n[287]), .ZN(R2_SB_n31) );
  INV_X1 R2_SB_U36 ( .A(R2_SB_n303), .ZN(R2_SB_n23) );
  INV_X1 R2_SB_U35 ( .A(R2_SB_n319), .ZN(R2_SB_n15) );
  INV_X1 R2_SB_U34 ( .A(R2_SB_n335), .ZN(R2_SB_n7) );
  INV_X1 R2_SB_U33 ( .A(R2_SB_n[286]), .ZN(R2_SB_n30) );
  INV_X1 R2_SB_U32 ( .A(R2_SB_n302), .ZN(R2_SB_n22) );
  INV_X1 R2_SB_U31 ( .A(R2_SB_n318), .ZN(R2_SB_n14) );
  INV_X1 R2_SB_U30 ( .A(R2_SB_n334), .ZN(R2_SB_n6) );
  INV_X1 R2_SB_U29 ( .A(R2_SB_n[282]), .ZN(R2_SB_n26) );
  INV_X1 R2_SB_U28 ( .A(R2_SB_n298), .ZN(R2_SB_n18) );
  INV_X1 R2_SB_U27 ( .A(R2_SB_n314), .ZN(R2_SB_n10) );
  INV_X1 R2_SB_U26 ( .A(R2_SB_n330), .ZN(R2_SB_n2) );
  INV_X1 R2_SB_U21 ( .A(R2_SB_n365), .ZN(R2_SB_n34) );
  BUF_X1 R2_SB_U20 ( .A(R2_SB_n363), .Z(R2_SB_n617) );
  BUF_X1 R2_SB_U18 ( .A(R2_SB_n361), .Z(R2_SB_n618) );
  NOR3_X1 R2_SB_U16 ( .A1(R2_SB_n617), .A2(R2_SB_n618), .A3(R2_SB_n616), .ZN(
        R2_SB_n373) );
  BUF_X1 R2_SB_U15 ( .A(R2_SB_n43), .Z(R2_SB_n621) );
  BUF_X1 R2_SB_U14 ( .A(R2_SB_n373), .Z(R2_SB_n615) );
  BUF_X1 R2_SB_U13 ( .A(R2_SB_n373), .Z(R2_SB_n614) );
  BUF_X1 R2_SB_U12 ( .A(R2_SB_n623), .Z(R2_SB_n624) );
  BUF_X1 R2_SB_U11 ( .A(R2_SB_n43), .Z(R2_SB_n622) );
  CLKBUF_X1 R2_SB_U9 ( .A(R2_SB_n619), .Z(R2_SB_n620) );
  CLKBUF_X1 R2_SB_U7 ( .A(R2_SB_n39), .Z(R2_SB_n625) );
  CLKBUF_X1 R2_SB_U6 ( .A(R2_SB_n39), .Z(R2_SB_n626) );
  NAND3_X1 R2_SB_U414 ( .A1(R2_SB_add_108_A_1_), .A2(R2_SB_n38), .A3(
        R2_SB_add_108_A_0_), .ZN(R2_SB_n423) );
  DLH_X1 R2_SB_ready_out_reg_39_ ( .G(R2_SB_n629), .D(R2_SB_n88), .Q(R2_n1555)
         );
  DFF_X1 R2_SB_temp_o_reg_39_ ( .D(R2_SB_n542), .CK(clk), .Q(R2_SB_n88) );
  DLH_X1 R2_SB_ready_out_reg_7_ ( .G(R2_SB_n629), .D(R2_SB_n56), .Q(R2_n1523)
         );
  DFF_X1 R2_SB_temp_o_reg_7_ ( .D(R2_SB_n541), .CK(clk), .Q(R2_SB_n56) );
  DLH_X1 R2_SB_ready_out_reg_71_ ( .G(R2_SB_n629), .D(R2_SB_n120), .Q(R2_n1587) );
  DFF_X1 R2_SB_temp_o_reg_71_ ( .D(R2_SB_n540), .CK(clk), .Q(R2_SB_n120) );
  DLH_X1 R2_SB_ready_out_reg_103_ ( .G(R2_SB_n629), .D(R2_SB_n152), .Q(
        R2_n1619) );
  DFF_X1 R2_SB_temp_o_reg_103_ ( .D(R2_SB_n539), .CK(clk), .Q(R2_SB_n152) );
  DLH_X1 R2_SB_ready_out_reg_38_ ( .G(R2_SB_n629), .D(R2_SB_n87), .Q(R2_n1554)
         );
  DFF_X1 R2_SB_temp_o_reg_38_ ( .D(R2_SB_n546), .CK(clk), .Q(R2_SB_n87) );
  DLH_X1 R2_SB_ready_out_reg_6_ ( .G(R2_SB_n628), .D(R2_SB_n55), .Q(R2_n1522)
         );
  DFF_X1 R2_SB_temp_o_reg_6_ ( .D(R2_SB_n545), .CK(clk), .Q(R2_SB_n55) );
  DLH_X1 R2_SB_ready_out_reg_70_ ( .G(R2_SB_n628), .D(R2_SB_n119), .Q(R2_n1586) );
  DFF_X1 R2_SB_temp_o_reg_70_ ( .D(R2_SB_n544), .CK(clk), .Q(R2_SB_n119) );
  DLH_X1 R2_SB_ready_out_reg_102_ ( .G(R2_SB_n628), .D(R2_SB_n151), .Q(
        R2_n1618) );
  DFF_X1 R2_SB_temp_o_reg_102_ ( .D(R2_SB_n543), .CK(clk), .Q(R2_SB_n151) );
  DLH_X1 R2_SB_ready_out_reg_37_ ( .G(R2_SB_n628), .D(R2_SB_n86), .Q(R2_n1553)
         );
  DFF_X1 R2_SB_temp_o_reg_37_ ( .D(R2_SB_n550), .CK(clk), .Q(R2_SB_n86) );
  DLH_X1 R2_SB_ready_out_reg_5_ ( .G(R2_SB_n628), .D(R2_SB_n54), .Q(R2_n1521)
         );
  DFF_X1 R2_SB_temp_o_reg_5_ ( .D(R2_SB_n549), .CK(clk), .Q(R2_SB_n54) );
  DLH_X1 R2_SB_ready_out_reg_69_ ( .G(R2_SB_n628), .D(R2_SB_n118), .Q(R2_n1585) );
  DFF_X1 R2_SB_temp_o_reg_69_ ( .D(R2_SB_n548), .CK(clk), .Q(R2_SB_n118) );
  DLH_X1 R2_SB_ready_out_reg_101_ ( .G(R2_SB_n628), .D(R2_SB_n150), .Q(
        R2_n1617) );
  DFF_X1 R2_SB_temp_o_reg_101_ ( .D(R2_SB_n547), .CK(clk), .Q(R2_SB_n150) );
  DLH_X1 R2_SB_ready_out_reg_36_ ( .G(R2_SB_n628), .D(R2_SB_n85), .Q(R2_n1552)
         );
  DFF_X1 R2_SB_temp_o_reg_36_ ( .D(R2_SB_n554), .CK(clk), .Q(R2_SB_n85) );
  DLH_X1 R2_SB_ready_out_reg_4_ ( .G(R2_SB_n628), .D(R2_SB_n53), .Q(R2_n1520)
         );
  DFF_X1 R2_SB_temp_o_reg_4_ ( .D(R2_SB_n553), .CK(clk), .Q(R2_SB_n53) );
  DLH_X1 R2_SB_ready_out_reg_68_ ( .G(R2_SB_n628), .D(R2_SB_n117), .Q(R2_n1584) );
  DFF_X1 R2_SB_temp_o_reg_68_ ( .D(R2_SB_n552), .CK(clk), .Q(R2_SB_n117) );
  DLH_X1 R2_SB_ready_out_reg_100_ ( .G(R2_SB_n628), .D(R2_SB_n149), .Q(
        R2_n1616) );
  DFF_X1 R2_SB_temp_o_reg_100_ ( .D(R2_SB_n551), .CK(clk), .Q(R2_SB_n149) );
  DLH_X1 R2_SB_ready_out_reg_35_ ( .G(R2_SB_n628), .D(R2_SB_n84), .Q(R2_n1551)
         );
  DFF_X1 R2_SB_temp_o_reg_35_ ( .D(R2_SB_n558), .CK(clk), .Q(R2_SB_n84) );
  DLH_X1 R2_SB_ready_out_reg_3_ ( .G(R2_SB_n628), .D(R2_SB_n52), .Q(R2_n1519)
         );
  DFF_X1 R2_SB_temp_o_reg_3_ ( .D(R2_SB_n557), .CK(clk), .Q(R2_SB_n52) );
  DLH_X1 R2_SB_ready_out_reg_67_ ( .G(R2_SB_n628), .D(R2_SB_n116), .Q(R2_n1583) );
  DFF_X1 R2_SB_temp_o_reg_67_ ( .D(R2_SB_n556), .CK(clk), .Q(R2_SB_n116) );
  DLH_X1 R2_SB_ready_out_reg_99_ ( .G(R2_SB_n628), .D(R2_SB_n148), .Q(R2_n1615) );
  DFF_X1 R2_SB_temp_o_reg_99_ ( .D(R2_SB_n555), .CK(clk), .Q(R2_SB_n148) );
  DLH_X1 R2_SB_ready_out_reg_34_ ( .G(R2_SB_n628), .D(R2_SB_n83), .Q(R2_n1550)
         );
  DFF_X1 R2_SB_temp_o_reg_34_ ( .D(R2_SB_n562), .CK(clk), .Q(R2_SB_n83) );
  DLH_X1 R2_SB_ready_out_reg_2_ ( .G(R2_SB_n628), .D(R2_SB_n51), .Q(R2_n1518)
         );
  DFF_X1 R2_SB_temp_o_reg_2_ ( .D(R2_SB_n561), .CK(clk), .Q(R2_SB_n51) );
  DLH_X1 R2_SB_ready_out_reg_66_ ( .G(R2_SB_n628), .D(R2_SB_n115), .Q(R2_n1582) );
  DFF_X1 R2_SB_temp_o_reg_66_ ( .D(R2_SB_n560), .CK(clk), .Q(R2_SB_n115) );
  DLH_X1 R2_SB_ready_out_reg_98_ ( .G(R2_SB_n628), .D(R2_SB_n147), .Q(R2_n1614) );
  DFF_X1 R2_SB_temp_o_reg_98_ ( .D(R2_SB_n559), .CK(clk), .Q(R2_SB_n147) );
  DLH_X1 R2_SB_ready_out_reg_33_ ( .G(R2_SB_n628), .D(R2_SB_n82), .Q(R2_n1549)
         );
  DFF_X1 R2_SB_temp_o_reg_33_ ( .D(R2_SB_n566), .CK(clk), .Q(R2_SB_n82) );
  DLH_X1 R2_SB_ready_out_reg_1_ ( .G(R2_SB_n628), .D(R2_SB_n50), .Q(R2_n1517)
         );
  DFF_X1 R2_SB_temp_o_reg_1_ ( .D(R2_SB_n565), .CK(clk), .Q(R2_SB_n50) );
  DLH_X1 R2_SB_ready_out_reg_65_ ( .G(R2_SB_n628), .D(R2_SB_n114), .Q(R2_n1581) );
  DFF_X1 R2_SB_temp_o_reg_65_ ( .D(R2_SB_n564), .CK(clk), .Q(R2_SB_n114) );
  DLH_X1 R2_SB_ready_out_reg_97_ ( .G(R2_SB_n628), .D(R2_SB_n146), .Q(R2_n1613) );
  DFF_X1 R2_SB_temp_o_reg_97_ ( .D(R2_SB_n563), .CK(clk), .Q(R2_SB_n146) );
  DLH_X1 R2_SB_ready_out_reg_32_ ( .G(R2_SB_n628), .D(R2_SB_n81), .Q(R2_n1548)
         );
  DFF_X1 R2_SB_temp_o_reg_32_ ( .D(R2_SB_n570), .CK(clk), .Q(R2_SB_n81) );
  DLH_X1 R2_SB_ready_out_reg_0_ ( .G(R2_SB_n628), .D(R2_SB_n49), .Q(R2_n1516)
         );
  DFF_X1 R2_SB_temp_o_reg_0_ ( .D(R2_SB_n569), .CK(clk), .Q(R2_SB_n49) );
  DLH_X1 R2_SB_ready_out_reg_64_ ( .G(R2_SB_n627), .D(R2_SB_n113), .Q(R2_n1580) );
  DFF_X1 R2_SB_temp_o_reg_64_ ( .D(R2_SB_n568), .CK(clk), .Q(R2_SB_n113) );
  DLH_X1 R2_SB_ready_out_reg_96_ ( .G(R2_SB_n627), .D(R2_SB_n145), .Q(R2_n1612) );
  DFF_X1 R2_SB_temp_o_reg_96_ ( .D(R2_SB_n567), .CK(clk), .Q(R2_SB_n145) );
  DLH_X1 R2_SB_sbox_s1_reg_0_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_0), .Q(
        R2_SB_n337) );
  DLH_X1 R2_SB_sbox_s1_reg_2_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_2), .Q(
        R2_SB_n339) );
  DLH_X1 R2_SB_sbox_s1_reg_3_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_3), .Q(
        R2_SB_n340) );
  DLH_X1 R2_SB_sbox_s1_reg_4_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_4), .Q(
        R2_SB_n341) );
  DLH_X1 R2_SB_sbox_s1_reg_5_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_5), .Q(
        R2_SB_n342) );
  DLH_X1 R2_SB_sbox_s1_reg_6_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_6), .Q(
        R2_SB_n343) );
  DLH_X1 R2_SB_sbox_s1_reg_7_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U10_Z_7), .Q(
        R2_SB_n344) );
  DLH_X1 R2_SB_ready_out_reg_47_ ( .G(R2_SB_n627), .D(R2_SB_n96), .Q(R2_n1563)
         );
  DFF_X1 R2_SB_temp_o_reg_47_ ( .D(R2_SB_n510), .CK(clk), .Q(R2_SB_n96) );
  DLH_X1 R2_SB_ready_out_reg_15_ ( .G(R2_SB_n627), .D(R2_SB_n64), .Q(R2_n1531)
         );
  DFF_X1 R2_SB_temp_o_reg_15_ ( .D(R2_SB_n509), .CK(clk), .Q(R2_SB_n64) );
  DLH_X1 R2_SB_ready_out_reg_79_ ( .G(R2_SB_n627), .D(R2_SB_n128), .Q(R2_n1595) );
  DFF_X1 R2_SB_temp_o_reg_79_ ( .D(R2_SB_n508), .CK(clk), .Q(R2_SB_n128) );
  DLH_X1 R2_SB_ready_out_reg_111_ ( .G(R2_SB_n627), .D(R2_SB_n160), .Q(
        R2_n1627) );
  DFF_X1 R2_SB_temp_o_reg_111_ ( .D(R2_SB_n507), .CK(clk), .Q(R2_SB_n160) );
  DLH_X1 R2_SB_ready_out_reg_46_ ( .G(R2_SB_n627), .D(R2_SB_n95), .Q(R2_n1562)
         );
  DFF_X1 R2_SB_temp_o_reg_46_ ( .D(R2_SB_n514), .CK(clk), .Q(R2_SB_n95) );
  DLH_X1 R2_SB_ready_out_reg_14_ ( .G(R2_SB_n627), .D(R2_SB_n63), .Q(R2_n1530)
         );
  DFF_X1 R2_SB_temp_o_reg_14_ ( .D(R2_SB_n513), .CK(clk), .Q(R2_SB_n63) );
  DLH_X1 R2_SB_ready_out_reg_78_ ( .G(R2_SB_n627), .D(R2_SB_n127), .Q(R2_n1594) );
  DFF_X1 R2_SB_temp_o_reg_78_ ( .D(R2_SB_n512), .CK(clk), .Q(R2_SB_n127) );
  DLH_X1 R2_SB_ready_out_reg_110_ ( .G(R2_SB_n627), .D(R2_SB_n159), .Q(
        R2_n1626) );
  DFF_X1 R2_SB_temp_o_reg_110_ ( .D(R2_SB_n511), .CK(clk), .Q(R2_SB_n159) );
  DLH_X1 R2_SB_ready_out_reg_45_ ( .G(R2_SB_n627), .D(R2_SB_n94), .Q(R2_n1561)
         );
  DFF_X1 R2_SB_temp_o_reg_45_ ( .D(R2_SB_n518), .CK(clk), .Q(R2_SB_n94) );
  DLH_X1 R2_SB_ready_out_reg_13_ ( .G(R2_SB_n627), .D(R2_SB_n62), .Q(R2_n1529)
         );
  DFF_X1 R2_SB_temp_o_reg_13_ ( .D(R2_SB_n517), .CK(clk), .Q(R2_SB_n62) );
  DLH_X1 R2_SB_ready_out_reg_77_ ( .G(R2_SB_n627), .D(R2_SB_n126), .Q(R2_n1593) );
  DFF_X1 R2_SB_temp_o_reg_77_ ( .D(R2_SB_n516), .CK(clk), .Q(R2_SB_n126) );
  DLH_X1 R2_SB_ready_out_reg_109_ ( .G(R2_SB_n627), .D(R2_SB_n158), .Q(
        R2_n1625) );
  DFF_X1 R2_SB_temp_o_reg_109_ ( .D(R2_SB_n515), .CK(clk), .Q(R2_SB_n158) );
  DLH_X1 R2_SB_ready_out_reg_44_ ( .G(R2_SB_n627), .D(R2_SB_n93), .Q(R2_n1560)
         );
  DFF_X1 R2_SB_temp_o_reg_44_ ( .D(R2_SB_n522), .CK(clk), .Q(R2_SB_n93) );
  DLH_X1 R2_SB_ready_out_reg_12_ ( .G(R2_SB_n627), .D(R2_SB_n61), .Q(R2_n1528)
         );
  DFF_X1 R2_SB_temp_o_reg_12_ ( .D(R2_SB_n521), .CK(clk), .Q(R2_SB_n61) );
  DLH_X1 R2_SB_ready_out_reg_76_ ( .G(R2_SB_n627), .D(R2_SB_n125), .Q(R2_n1592) );
  DFF_X1 R2_SB_temp_o_reg_76_ ( .D(R2_SB_n520), .CK(clk), .Q(R2_SB_n125) );
  DLH_X1 R2_SB_ready_out_reg_108_ ( .G(R2_SB_n627), .D(R2_SB_n157), .Q(
        R2_n1624) );
  DFF_X1 R2_SB_temp_o_reg_108_ ( .D(R2_SB_n519), .CK(clk), .Q(R2_SB_n157) );
  DLH_X1 R2_SB_ready_out_reg_43_ ( .G(R2_SB_n627), .D(R2_SB_n92), .Q(R2_n1559)
         );
  DFF_X1 R2_SB_temp_o_reg_43_ ( .D(R2_SB_n526), .CK(clk), .Q(R2_SB_n92) );
  DLH_X1 R2_SB_ready_out_reg_11_ ( .G(R2_SB_n627), .D(R2_SB_n60), .Q(R2_n1527)
         );
  DFF_X1 R2_SB_temp_o_reg_11_ ( .D(R2_SB_n525), .CK(clk), .Q(R2_SB_n60) );
  DLH_X1 R2_SB_ready_out_reg_75_ ( .G(R2_SB_n627), .D(R2_SB_n124), .Q(R2_n1591) );
  DFF_X1 R2_SB_temp_o_reg_75_ ( .D(R2_SB_n524), .CK(clk), .Q(R2_SB_n124) );
  DLH_X1 R2_SB_ready_out_reg_107_ ( .G(R2_SB_n627), .D(R2_SB_n156), .Q(
        R2_n1623) );
  DFF_X1 R2_SB_temp_o_reg_107_ ( .D(R2_SB_n523), .CK(clk), .Q(R2_SB_n156) );
  DLH_X1 R2_SB_ready_out_reg_42_ ( .G(R2_SB_n627), .D(R2_SB_n91), .Q(R2_n1558)
         );
  DFF_X1 R2_SB_temp_o_reg_42_ ( .D(R2_SB_n530), .CK(clk), .Q(R2_SB_n91) );
  DLH_X1 R2_SB_ready_out_reg_10_ ( .G(R2_SB_n627), .D(R2_SB_n59), .Q(R2_n1526)
         );
  DFF_X1 R2_SB_temp_o_reg_10_ ( .D(R2_SB_n529), .CK(clk), .Q(R2_SB_n59) );
  DLH_X1 R2_SB_ready_out_reg_74_ ( .G(R2_SB_n627), .D(R2_SB_n123), .Q(R2_n1590) );
  DFF_X1 R2_SB_temp_o_reg_74_ ( .D(R2_SB_n528), .CK(clk), .Q(R2_SB_n123) );
  DLH_X1 R2_SB_ready_out_reg_106_ ( .G(R2_SB_n276), .D(R2_SB_n155), .Q(
        R2_n1622) );
  DFF_X1 R2_SB_temp_o_reg_106_ ( .D(R2_SB_n527), .CK(clk), .Q(R2_SB_n155) );
  DLH_X1 R2_SB_ready_out_reg_41_ ( .G(R2_SB_n276), .D(R2_SB_n90), .Q(R2_n1557)
         );
  DFF_X1 R2_SB_temp_o_reg_41_ ( .D(R2_SB_n534), .CK(clk), .Q(R2_SB_n90) );
  DLH_X1 R2_SB_ready_out_reg_9_ ( .G(R2_SB_n276), .D(R2_SB_n58), .Q(R2_n1525)
         );
  DFF_X1 R2_SB_temp_o_reg_9_ ( .D(R2_SB_n533), .CK(clk), .Q(R2_SB_n58) );
  DLH_X1 R2_SB_ready_out_reg_73_ ( .G(R2_SB_n276), .D(R2_SB_n122), .Q(R2_n1589) );
  DFF_X1 R2_SB_temp_o_reg_73_ ( .D(R2_SB_n532), .CK(clk), .Q(R2_SB_n122) );
  DLH_X1 R2_SB_ready_out_reg_105_ ( .G(R2_SB_n276), .D(R2_SB_n154), .Q(
        R2_n1621) );
  DFF_X1 R2_SB_temp_o_reg_105_ ( .D(R2_SB_n531), .CK(clk), .Q(R2_SB_n154) );
  DLH_X1 R2_SB_ready_out_reg_40_ ( .G(R2_SB_n276), .D(R2_SB_n89), .Q(R2_n1556)
         );
  DFF_X1 R2_SB_temp_o_reg_40_ ( .D(R2_SB_n538), .CK(clk), .Q(R2_SB_n89) );
  DLH_X1 R2_SB_ready_out_reg_8_ ( .G(R2_SB_n276), .D(R2_SB_n57), .Q(R2_n1524)
         );
  DFF_X1 R2_SB_temp_o_reg_8_ ( .D(R2_SB_n537), .CK(clk), .Q(R2_SB_n57) );
  DLH_X1 R2_SB_ready_out_reg_72_ ( .G(R2_SB_n276), .D(R2_SB_n121), .Q(R2_n1588) );
  DFF_X1 R2_SB_temp_o_reg_72_ ( .D(R2_SB_n536), .CK(clk), .Q(R2_SB_n121) );
  DLH_X1 R2_SB_ready_out_reg_104_ ( .G(R2_SB_n276), .D(R2_SB_n153), .Q(
        R2_n1620) );
  DFF_X1 R2_SB_temp_o_reg_104_ ( .D(R2_SB_n535), .CK(clk), .Q(R2_SB_n153) );
  DLH_X1 R2_SB_sbox_s2_reg_0_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_0), .Q(
        R2_SB_n321) );
  DLH_X1 R2_SB_sbox_s2_reg_2_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_2), .Q(
        R2_SB_n323) );
  DLH_X1 R2_SB_sbox_s2_reg_3_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_3), .Q(
        R2_SB_n324) );
  DLH_X1 R2_SB_sbox_s2_reg_4_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_4), .Q(
        R2_SB_n325) );
  DLH_X1 R2_SB_sbox_s2_reg_5_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_5), .Q(
        R2_SB_n326) );
  DLH_X1 R2_SB_sbox_s2_reg_6_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_6), .Q(
        R2_SB_n327) );
  DLH_X1 R2_SB_sbox_s2_reg_7_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U9_Z_7), .Q(
        R2_SB_n328) );
  DLH_X1 R2_SB_ready_out_reg_55_ ( .G(R2_SB_n276), .D(R2_SB_n104), .Q(R2_n1571) );
  DFF_X1 R2_SB_temp_o_reg_55_ ( .D(R2_SB_n478), .CK(clk), .Q(R2_SB_n104) );
  DLH_X1 R2_SB_ready_out_reg_23_ ( .G(R2_SB_n276), .D(R2_SB_n72), .Q(R2_n1539)
         );
  DFF_X1 R2_SB_temp_o_reg_23_ ( .D(R2_SB_n477), .CK(clk), .Q(R2_SB_n72) );
  DLH_X1 R2_SB_ready_out_reg_87_ ( .G(R2_SB_n276), .D(R2_SB_n136), .Q(R2_n1603) );
  DFF_X1 R2_SB_temp_o_reg_87_ ( .D(R2_SB_n476), .CK(clk), .Q(R2_SB_n136) );
  DLH_X1 R2_SB_ready_out_reg_119_ ( .G(R2_SB_n276), .D(R2_SB_n168), .Q(
        R2_n1635) );
  DFF_X1 R2_SB_temp_o_reg_119_ ( .D(R2_SB_n475), .CK(clk), .Q(R2_SB_n168) );
  DLH_X1 R2_SB_ready_out_reg_54_ ( .G(R2_SB_n276), .D(R2_SB_n103), .Q(R2_n1570) );
  DFF_X1 R2_SB_temp_o_reg_54_ ( .D(R2_SB_n482), .CK(clk), .Q(R2_SB_n103) );
  DLH_X1 R2_SB_ready_out_reg_22_ ( .G(R2_SB_n276), .D(R2_SB_n71), .Q(R2_n1538)
         );
  DFF_X1 R2_SB_temp_o_reg_22_ ( .D(R2_SB_n481), .CK(clk), .Q(R2_SB_n71) );
  DLH_X1 R2_SB_ready_out_reg_86_ ( .G(R2_SB_n276), .D(R2_SB_n135), .Q(R2_n1602) );
  DFF_X1 R2_SB_temp_o_reg_86_ ( .D(R2_SB_n480), .CK(clk), .Q(R2_SB_n135) );
  DLH_X1 R2_SB_ready_out_reg_118_ ( .G(R2_SB_n276), .D(R2_SB_n167), .Q(
        R2_n1634) );
  DFF_X1 R2_SB_temp_o_reg_118_ ( .D(R2_SB_n479), .CK(clk), .Q(R2_SB_n167) );
  DLH_X1 R2_SB_ready_out_reg_53_ ( .G(R2_SB_n276), .D(R2_SB_n102), .Q(R2_n1569) );
  DFF_X1 R2_SB_temp_o_reg_53_ ( .D(R2_SB_n486), .CK(clk), .Q(R2_SB_n102) );
  DLH_X1 R2_SB_ready_out_reg_21_ ( .G(R2_SB_n276), .D(R2_SB_n70), .Q(R2_n1537)
         );
  DFF_X1 R2_SB_temp_o_reg_21_ ( .D(R2_SB_n485), .CK(clk), .Q(R2_SB_n70) );
  DLH_X1 R2_SB_ready_out_reg_85_ ( .G(R2_SB_n276), .D(R2_SB_n134), .Q(R2_n1601) );
  DFF_X1 R2_SB_temp_o_reg_85_ ( .D(R2_SB_n484), .CK(clk), .Q(R2_SB_n134) );
  DLH_X1 R2_SB_ready_out_reg_117_ ( .G(R2_SB_n276), .D(R2_SB_n166), .Q(
        R2_n1633) );
  DFF_X1 R2_SB_temp_o_reg_117_ ( .D(R2_SB_n483), .CK(clk), .Q(R2_SB_n166) );
  DLH_X1 R2_SB_ready_out_reg_52_ ( .G(R2_SB_n276), .D(R2_SB_n101), .Q(R2_n1568) );
  DFF_X1 R2_SB_temp_o_reg_52_ ( .D(R2_SB_n490), .CK(clk), .Q(R2_SB_n101) );
  DLH_X1 R2_SB_ready_out_reg_20_ ( .G(R2_SB_n276), .D(R2_SB_n69), .Q(R2_n1536)
         );
  DFF_X1 R2_SB_temp_o_reg_20_ ( .D(R2_SB_n489), .CK(clk), .Q(R2_SB_n69) );
  DLH_X1 R2_SB_ready_out_reg_84_ ( .G(R2_SB_n276), .D(R2_SB_n133), .Q(R2_n1600) );
  DFF_X1 R2_SB_temp_o_reg_84_ ( .D(R2_SB_n488), .CK(clk), .Q(R2_SB_n133) );
  DLH_X1 R2_SB_ready_out_reg_116_ ( .G(R2_SB_n276), .D(R2_SB_n165), .Q(
        R2_n1632) );
  DFF_X1 R2_SB_temp_o_reg_116_ ( .D(R2_SB_n487), .CK(clk), .Q(R2_SB_n165) );
  DLH_X1 R2_SB_ready_out_reg_51_ ( .G(R2_SB_n629), .D(R2_SB_n100), .Q(R2_n1567) );
  DFF_X1 R2_SB_temp_o_reg_51_ ( .D(R2_SB_n494), .CK(clk), .Q(R2_SB_n100) );
  DLH_X1 R2_SB_ready_out_reg_19_ ( .G(R2_SB_n629), .D(R2_SB_n68), .Q(R2_n1535)
         );
  DFF_X1 R2_SB_temp_o_reg_19_ ( .D(R2_SB_n493), .CK(clk), .Q(R2_SB_n68) );
  DLH_X1 R2_SB_ready_out_reg_83_ ( .G(R2_SB_n629), .D(R2_SB_n132), .Q(R2_n1599) );
  DFF_X1 R2_SB_temp_o_reg_83_ ( .D(R2_SB_n492), .CK(clk), .Q(R2_SB_n132) );
  DLH_X1 R2_SB_ready_out_reg_115_ ( .G(R2_SB_n629), .D(R2_SB_n164), .Q(
        R2_n1631) );
  DFF_X1 R2_SB_temp_o_reg_115_ ( .D(R2_SB_n491), .CK(clk), .Q(R2_SB_n164) );
  DLH_X1 R2_SB_ready_out_reg_50_ ( .G(R2_SB_n629), .D(R2_SB_n99), .Q(R2_n1566)
         );
  DFF_X1 R2_SB_temp_o_reg_50_ ( .D(R2_SB_n498), .CK(clk), .Q(R2_SB_n99) );
  DLH_X1 R2_SB_ready_out_reg_18_ ( .G(R2_SB_n629), .D(R2_SB_n67), .Q(R2_n1534)
         );
  DFF_X1 R2_SB_temp_o_reg_18_ ( .D(R2_SB_n497), .CK(clk), .Q(R2_SB_n67) );
  DLH_X1 R2_SB_ready_out_reg_82_ ( .G(R2_SB_n629), .D(R2_SB_n131), .Q(R2_n1598) );
  DFF_X1 R2_SB_temp_o_reg_82_ ( .D(R2_SB_n496), .CK(clk), .Q(R2_SB_n131) );
  DLH_X1 R2_SB_ready_out_reg_114_ ( .G(R2_SB_n629), .D(R2_SB_n163), .Q(
        R2_n1630) );
  DFF_X1 R2_SB_temp_o_reg_114_ ( .D(R2_SB_n495), .CK(clk), .Q(R2_SB_n163) );
  DLH_X1 R2_SB_ready_out_reg_49_ ( .G(R2_SB_n629), .D(R2_SB_n98), .Q(R2_n1565)
         );
  DFF_X1 R2_SB_temp_o_reg_49_ ( .D(R2_SB_n502), .CK(clk), .Q(R2_SB_n98) );
  DLH_X1 R2_SB_ready_out_reg_17_ ( .G(R2_SB_n629), .D(R2_SB_n66), .Q(R2_n1533)
         );
  DFF_X1 R2_SB_temp_o_reg_17_ ( .D(R2_SB_n501), .CK(clk), .Q(R2_SB_n66) );
  DLH_X1 R2_SB_ready_out_reg_81_ ( .G(R2_SB_n629), .D(R2_SB_n130), .Q(R2_n1597) );
  DFF_X1 R2_SB_temp_o_reg_81_ ( .D(R2_SB_n500), .CK(clk), .Q(R2_SB_n130) );
  DLH_X1 R2_SB_ready_out_reg_113_ ( .G(R2_SB_n629), .D(R2_SB_n162), .Q(
        R2_n1629) );
  DFF_X1 R2_SB_temp_o_reg_113_ ( .D(R2_SB_n499), .CK(clk), .Q(R2_SB_n162) );
  DLH_X1 R2_SB_ready_out_reg_48_ ( .G(R2_SB_n629), .D(R2_SB_n97), .Q(R2_n1564)
         );
  DFF_X1 R2_SB_temp_o_reg_48_ ( .D(R2_SB_n506), .CK(clk), .Q(R2_SB_n97) );
  DLH_X1 R2_SB_ready_out_reg_16_ ( .G(R2_SB_n629), .D(R2_SB_n65), .Q(R2_n1532)
         );
  DFF_X1 R2_SB_temp_o_reg_16_ ( .D(R2_SB_n505), .CK(clk), .Q(R2_SB_n65) );
  DLH_X1 R2_SB_ready_out_reg_80_ ( .G(R2_SB_n629), .D(R2_SB_n129), .Q(R2_n1596) );
  DFF_X1 R2_SB_temp_o_reg_80_ ( .D(R2_SB_n504), .CK(clk), .Q(R2_SB_n129) );
  DLH_X1 R2_SB_ready_out_reg_112_ ( .G(R2_SB_n629), .D(R2_SB_n161), .Q(
        R2_n1628) );
  DFF_X1 R2_SB_temp_o_reg_112_ ( .D(R2_SB_n503), .CK(clk), .Q(R2_SB_n161) );
  DLH_X1 R2_SB_sbox_s3_reg_0_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_0), .Q(
        R2_SB_n305) );
  DLH_X1 R2_SB_sbox_s3_reg_2_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_2), .Q(
        R2_SB_n307) );
  DLH_X1 R2_SB_sbox_s3_reg_3_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_3), .Q(
        R2_SB_n308) );
  DLH_X1 R2_SB_sbox_s3_reg_4_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_4), .Q(
        R2_SB_n309) );
  DLH_X1 R2_SB_sbox_s3_reg_5_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_5), .Q(
        R2_SB_n310) );
  DLH_X1 R2_SB_sbox_s3_reg_6_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_6), .Q(
        R2_SB_n311) );
  DLH_X1 R2_SB_sbox_s3_reg_7_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U8_Z_7), .Q(
        R2_SB_n312) );
  DLH_X1 R2_SB_ready_out_reg_63_ ( .G(R2_SB_n276), .D(R2_SB_n112), .Q(R2_n1579) );
  DFF_X1 R2_SB_temp_o_reg_63_ ( .D(R2_SB_n446), .CK(clk), .Q(R2_SB_n112) );
  DLH_X1 R2_SB_ready_out_reg_31_ ( .G(R2_SB_n629), .D(R2_SB_n80), .Q(R2_n1547)
         );
  DFF_X1 R2_SB_temp_o_reg_31_ ( .D(R2_SB_n445), .CK(clk), .Q(R2_SB_n80) );
  DLH_X1 R2_SB_ready_out_reg_95_ ( .G(R2_SB_n628), .D(R2_SB_n144), .Q(R2_n1611) );
  DFF_X1 R2_SB_temp_o_reg_95_ ( .D(R2_SB_n444), .CK(clk), .Q(R2_SB_n144) );
  DLH_X1 R2_SB_ready_out_reg_127_ ( .G(R2_SB_n629), .D(R2_SB_n176), .Q(
        R2_n1643) );
  DFF_X1 R2_SB_temp_o_reg_127_ ( .D(R2_SB_n443), .CK(clk), .Q(R2_SB_n176) );
  DLH_X1 R2_SB_ready_out_reg_62_ ( .G(R2_SB_n629), .D(R2_SB_n111), .Q(R2_n1578) );
  DFF_X1 R2_SB_temp_o_reg_62_ ( .D(R2_SB_n450), .CK(clk), .Q(R2_SB_n111) );
  DLH_X1 R2_SB_ready_out_reg_30_ ( .G(R2_SB_n629), .D(R2_SB_n79), .Q(R2_n1546)
         );
  DFF_X1 R2_SB_temp_o_reg_30_ ( .D(R2_SB_n449), .CK(clk), .Q(R2_SB_n79) );
  DLH_X1 R2_SB_ready_out_reg_94_ ( .G(R2_SB_n629), .D(R2_SB_n143), .Q(R2_n1610) );
  DFF_X1 R2_SB_temp_o_reg_94_ ( .D(R2_SB_n448), .CK(clk), .Q(R2_SB_n143) );
  DLH_X1 R2_SB_ready_out_reg_126_ ( .G(R2_SB_n629), .D(R2_SB_n175), .Q(
        R2_n1642) );
  DFF_X1 R2_SB_temp_o_reg_126_ ( .D(R2_SB_n447), .CK(clk), .Q(R2_SB_n175) );
  DLH_X1 R2_SB_ready_out_reg_61_ ( .G(R2_SB_n628), .D(R2_SB_n110), .Q(R2_n1577) );
  DFF_X1 R2_SB_temp_o_reg_61_ ( .D(R2_SB_n454), .CK(clk), .Q(R2_SB_n110) );
  DLH_X1 R2_SB_ready_out_reg_29_ ( .G(R2_SB_n627), .D(R2_SB_n78), .Q(R2_n1545)
         );
  DFF_X1 R2_SB_temp_o_reg_29_ ( .D(R2_SB_n453), .CK(clk), .Q(R2_SB_n78) );
  DLH_X1 R2_SB_ready_out_reg_93_ ( .G(R2_SB_n629), .D(R2_SB_n142), .Q(R2_n1609) );
  DFF_X1 R2_SB_temp_o_reg_93_ ( .D(R2_SB_n452), .CK(clk), .Q(R2_SB_n142) );
  DLH_X1 R2_SB_ready_out_reg_125_ ( .G(R2_SB_n628), .D(R2_SB_n174), .Q(
        R2_n1641) );
  DFF_X1 R2_SB_temp_o_reg_125_ ( .D(R2_SB_n451), .CK(clk), .Q(R2_SB_n174) );
  DLH_X1 R2_SB_ready_out_reg_60_ ( .G(R2_SB_n627), .D(R2_SB_n109), .Q(R2_n1576) );
  DFF_X1 R2_SB_temp_o_reg_60_ ( .D(R2_SB_n458), .CK(clk), .Q(R2_SB_n109) );
  DLH_X1 R2_SB_ready_out_reg_28_ ( .G(R2_SB_n629), .D(R2_SB_n77), .Q(R2_n1544)
         );
  DFF_X1 R2_SB_temp_o_reg_28_ ( .D(R2_SB_n457), .CK(clk), .Q(R2_SB_n77) );
  DLH_X1 R2_SB_ready_out_reg_92_ ( .G(R2_SB_n628), .D(R2_SB_n141), .Q(R2_n1608) );
  DFF_X1 R2_SB_temp_o_reg_92_ ( .D(R2_SB_n456), .CK(clk), .Q(R2_SB_n141) );
  DLH_X1 R2_SB_ready_out_reg_124_ ( .G(R2_SB_n627), .D(R2_SB_n173), .Q(
        R2_n1640) );
  DFF_X1 R2_SB_temp_o_reg_124_ ( .D(R2_SB_n455), .CK(clk), .Q(R2_SB_n173) );
  DLH_X1 R2_SB_ready_out_reg_59_ ( .G(R2_SB_n628), .D(R2_SB_n108), .Q(R2_n1575) );
  DFF_X1 R2_SB_temp_o_reg_59_ ( .D(R2_SB_n462), .CK(clk), .Q(R2_SB_n108) );
  DLH_X1 R2_SB_ready_out_reg_27_ ( .G(R2_SB_n627), .D(R2_SB_n76), .Q(R2_n1543)
         );
  DFF_X1 R2_SB_temp_o_reg_27_ ( .D(R2_SB_n461), .CK(clk), .Q(R2_SB_n76) );
  DLH_X1 R2_SB_ready_out_reg_91_ ( .G(R2_SB_n629), .D(R2_SB_n140), .Q(R2_n1607) );
  DFF_X1 R2_SB_temp_o_reg_91_ ( .D(R2_SB_n460), .CK(clk), .Q(R2_SB_n140) );
  DLH_X1 R2_SB_ready_out_reg_123_ ( .G(R2_SB_n628), .D(R2_SB_n172), .Q(
        R2_n1639) );
  DFF_X1 R2_SB_temp_o_reg_123_ ( .D(R2_SB_n459), .CK(clk), .Q(R2_SB_n172) );
  DLH_X1 R2_SB_ready_out_reg_58_ ( .G(R2_SB_n276), .D(R2_SB_n107), .Q(R2_n1574) );
  DFF_X1 R2_SB_temp_o_reg_58_ ( .D(R2_SB_n466), .CK(clk), .Q(R2_SB_n107) );
  DLH_X1 R2_SB_ready_out_reg_26_ ( .G(R2_SB_n276), .D(R2_SB_n75), .Q(R2_n1542)
         );
  DFF_X1 R2_SB_temp_o_reg_26_ ( .D(R2_SB_n465), .CK(clk), .Q(R2_SB_n75) );
  DLH_X1 R2_SB_ready_out_reg_90_ ( .G(R2_SB_n276), .D(R2_SB_n139), .Q(R2_n1606) );
  DFF_X1 R2_SB_temp_o_reg_90_ ( .D(R2_SB_n464), .CK(clk), .Q(R2_SB_n139) );
  DLH_X1 R2_SB_ready_out_reg_122_ ( .G(R2_SB_n628), .D(R2_SB_n171), .Q(
        R2_n1638) );
  DFF_X1 R2_SB_temp_o_reg_122_ ( .D(R2_SB_n463), .CK(clk), .Q(R2_SB_n171) );
  DLH_X1 R2_SB_ready_out_reg_57_ ( .G(R2_SB_n629), .D(R2_SB_n106), .Q(R2_n1573) );
  DFF_X1 R2_SB_temp_o_reg_57_ ( .D(R2_SB_n470), .CK(clk), .Q(R2_SB_n106) );
  DLH_X1 R2_SB_ready_out_reg_25_ ( .G(R2_SB_n628), .D(R2_SB_n74), .Q(R2_n1541)
         );
  DFF_X1 R2_SB_temp_o_reg_25_ ( .D(R2_SB_n469), .CK(clk), .Q(R2_SB_n74) );
  DLH_X1 R2_SB_ready_out_reg_89_ ( .G(R2_SB_n627), .D(R2_SB_n138), .Q(R2_n1605) );
  DFF_X1 R2_SB_temp_o_reg_89_ ( .D(R2_SB_n468), .CK(clk), .Q(R2_SB_n138) );
  DLH_X1 R2_SB_ready_out_reg_121_ ( .G(R2_SB_n629), .D(R2_SB_n170), .Q(
        R2_n1637) );
  DFF_X1 R2_SB_temp_o_reg_121_ ( .D(R2_SB_n467), .CK(clk), .Q(R2_SB_n170) );
  DLH_X1 R2_SB_ready_out_reg_56_ ( .G(R2_SB_n627), .D(R2_SB_n105), .Q(R2_n1572) );
  DFF_X1 R2_SB_temp_o_reg_56_ ( .D(R2_SB_n474), .CK(clk), .Q(R2_SB_n105) );
  DLH_X1 R2_SB_ready_out_reg_24_ ( .G(R2_SB_n627), .D(R2_SB_n73), .Q(R2_n1540)
         );
  DFF_X1 R2_SB_temp_o_reg_24_ ( .D(R2_SB_n473), .CK(clk), .Q(R2_SB_n73) );
  DLH_X1 R2_SB_ready_out_reg_88_ ( .G(R2_SB_n627), .D(R2_SB_n137), .Q(R2_n1604) );
  DFF_X1 R2_SB_temp_o_reg_88_ ( .D(R2_SB_n472), .CK(clk), .Q(R2_SB_n137) );
  DLH_X1 R2_SB_ready_out_reg_120_ ( .G(R2_SB_n629), .D(R2_SB_n169), .Q(
        R2_n1636) );
  DFF_X1 R2_SB_temp_o_reg_120_ ( .D(R2_SB_n471), .CK(clk), .Q(R2_SB_n169) );
  DLH_X1 R2_SB_sbox_s4_reg_0_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_0), .Q(
        R2_SB_n289) );
  DLH_X1 R2_SB_sbox_s4_reg_2_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_2), .Q(
        R2_SB_n291) );
  DLH_X1 R2_SB_sbox_s4_reg_3_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_3), .Q(
        R2_SB_n292) );
  DLH_X1 R2_SB_sbox_s4_reg_4_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_4), .Q(
        R2_SB_n293) );
  DLH_X1 R2_SB_sbox_s4_reg_5_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_5), .Q(
        R2_SB_n294) );
  DLH_X1 R2_SB_sbox_s4_reg_6_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_6), .Q(
        R2_SB_n295) );
  DLH_X1 R2_SB_sbox_s4_reg_7_ ( .G(R2_SB_U11_Z_0), .D(R2_SB_U7_Z_7), .Q(
        R2_SB_n296) );
  DFF_X1 R2_SB_ready_reg ( .D(R2_SB_n572), .CK(clk), .Q(R2_n1515) );
  DFF_X1 R2_SB_cnt_reg_3_ ( .D(R2_SB_n33), .CK(clk), .Q(R2_SB_add_108_A_3_) );
  DFF_X1 R2_SB_cnt_reg_2_ ( .D(R2_SB_U4_Z_2), .CK(clk), .Q(R2_SB_add_108_A_2_), 
        .QN(R2_SB_n35) );
  DFF_X1 R2_SB_cnt_reg_1_ ( .D(R2_SB_U4_Z_1), .CK(clk), .Q(R2_SB_add_108_A_1_), 
        .QN(R2_SB_n36) );
  DFF_X1 R2_SB_cnt_reg_0_ ( .D(R2_SB_U4_Z_0), .CK(clk), .Q(R2_SB_add_108_A_0_), 
        .QN(R2_SB_n37) );
  INV_X1 R2_SB_SB1_U466 ( .A(R2_SB_SB1_n453), .ZN(R2_SB_SB1_n452) );
  INV_X1 R2_SB_SB1_U465 ( .A(R2_SB_n338), .ZN(R2_SB_SB1_n89) );
  INV_X1 R2_SB_SB1_U419 ( .A(R2_SB_n337), .ZN(R2_SB_SB1_n453) );
  NAND2_X1 R2_SB_SB1_U418 ( .A1(R2_SB_n338), .A2(R2_SB_n343), .ZN(
        R2_SB_SB1_n705) );
  AOI22_X1 R2_SB_SB1_U417 ( .A1(R2_SB_SB1_n779), .A2(R2_SB_SB1_n760), .B1(
        R2_SB_SB1_n877), .B2(R2_SB_SB1_n792), .ZN(R2_SB_SB1_n761) );
  OAI21_X1 R2_SB_SB1_U416 ( .B1(R2_SB_SB1_n759), .B2(R2_SB_SB1_n900), .A(
        R2_SB_SB1_n758), .ZN(R2_SB_SB1_n763) );
  AOI222_X1 R2_SB_SB1_U415 ( .A1(R2_SB_SB1_n742), .A2(R2_SB_n342), .B1(
        R2_SB_SB1_n778), .B2(R2_SB_SB1_n748), .C1(R2_SB_SB1_n747), .C2(
        R2_SB_SB1_n656), .ZN(R2_SB_SB1_n657) );
  NAND2_X1 R2_SB_SB1_U414 ( .A1(R2_SB_SB1_n743), .A2(R2_SB_n344), .ZN(
        R2_SB_SB1_n472) );
  AOI21_X1 R2_SB_SB1_U413 ( .B1(R2_SB_SB1_n835), .B2(R2_SB_SB1_n837), .A(
        R2_SB_SB1_n859), .ZN(R2_SB_SB1_n474) );
  OAI21_X1 R2_SB_SB1_U412 ( .B1(R2_SB_SB1_n474), .B2(R2_SB_SB1_n473), .A(
        R2_SB_SB1_n813), .ZN(R2_SB_SB1_n475) );
  OAI22_X1 R2_SB_SB1_U411 ( .A1(R2_SB_SB1_n829), .A2(R2_SB_SB1_n847), .B1(
        R2_SB_SB1_n845), .B2(R2_SB_SB1_n826), .ZN(R2_SB_SB1_n714) );
  NOR2_X1 R2_SB_SB1_U410 ( .A1(R2_SB_n344), .A2(R2_SB_SB1_n863), .ZN(
        R2_SB_SB1_n535) );
  OAI21_X1 R2_SB_SB1_U409 ( .B1(R2_SB_SB1_n855), .B2(R2_SB_SB1_n829), .A(
        R2_SB_SB1_n745), .ZN(R2_SB_SB1_n746) );
  AOI221_X1 R2_SB_SB1_U408 ( .B1(R2_SB_SB1_n805), .B2(R2_SB_SB1_n748), .C1(
        R2_SB_SB1_n747), .C2(R2_SB_SB1_n780), .A(R2_SB_SB1_n746), .ZN(
        R2_SB_SB1_n749) );
  AOI22_X1 R2_SB_SB1_U407 ( .A1(R2_SB_SB1_n742), .A2(R2_SB_n342), .B1(
        R2_SB_SB1_n778), .B2(R2_SB_SB1_n771), .ZN(R2_SB_SB1_n750) );
  OAI211_X1 R2_SB_SB1_U406 ( .C1(R2_SB_SB1_n828), .C2(R2_SB_SB1_n847), .A(
        R2_SB_SB1_n750), .B(R2_SB_SB1_n749), .ZN(R2_SB_SB1_n751) );
  NOR2_X1 R2_SB_SB1_U405 ( .A1(R2_SB_n342), .A2(R2_SB_SB1_n830), .ZN(
        R2_SB_SB1_n724) );
  NOR2_X1 R2_SB_SB1_U404 ( .A1(R2_SB_SB1_n826), .A2(R2_SB_n340), .ZN(
        R2_SB_SB1_n463) );
  OAI22_X1 R2_SB_SB1_U403 ( .A1(R2_SB_n344), .A2(R2_SB_SB1_n876), .B1(
        R2_SB_SB1_n858), .B2(R2_SB_SB1_n901), .ZN(R2_SB_SB1_n760) );
  NOR3_X1 R2_SB_SB1_U402 ( .A1(R2_SB_SB1_n890), .A2(R2_SB_n342), .A3(
        R2_SB_n338), .ZN(R2_SB_SB1_n613) );
  OAI22_X1 R2_SB_SB1_U401 ( .A1(R2_SB_SB1_n89), .A2(R2_SB_SB1_n898), .B1(
        R2_SB_SB1_n628), .B2(R2_SB_SB1_n907), .ZN(R2_SB_SB1_n614) );
  NOR3_X1 R2_SB_SB1_U400 ( .A1(R2_SB_SB1_n614), .A2(R2_SB_SB1_n722), .A3(
        R2_SB_SB1_n613), .ZN(R2_SB_SB1_n623) );
  NOR3_X1 R2_SB_SB1_U399 ( .A1(R2_SB_SB1_n863), .A2(R2_SB_n344), .A3(
        R2_SB_SB1_n814), .ZN(R2_SB_SB1_n797) );
  AOI22_X1 R2_SB_SB1_U398 ( .A1(R2_SB_SB1_n628), .A2(R2_SB_SB1_n627), .B1(
        R2_SB_n339), .B2(R2_SB_SB1_n730), .ZN(R2_SB_SB1_n630) );
  OAI222_X1 R2_SB_SB1_U397 ( .A1(R2_SB_SB1_n837), .A2(R2_SB_SB1_n573), .B1(
        R2_SB_n337), .B2(R2_SB_SB1_n468), .C1(R2_SB_n338), .C2(R2_SB_SB1_n677), 
        .ZN(R2_SB_SB1_n483) );
  OAI221_X1 R2_SB_SB1_U396 ( .B1(R2_SB_n340), .B2(R2_SB_SB1_n581), .C1(
        R2_SB_SB1_n476), .C2(R2_SB_SB1_n878), .A(R2_SB_SB1_n475), .ZN(
        R2_SB_SB1_n482) );
  OAI22_X1 R2_SB_SB1_U395 ( .A1(R2_SB_SB1_n840), .A2(R2_SB_SB1_n800), .B1(
        R2_SB_SB1_n480), .B2(R2_SB_SB1_n453), .ZN(R2_SB_SB1_n481) );
  NOR4_X1 R2_SB_SB1_U394 ( .A1(R2_SB_SB1_n484), .A2(R2_SB_SB1_n483), .A3(
        R2_SB_SB1_n482), .A4(R2_SB_SB1_n481), .ZN(R2_SB_SB1_n485) );
  NOR2_X1 R2_SB_SB1_U393 ( .A1(R2_SB_SB1_n868), .A2(R2_SB_n344), .ZN(
        R2_SB_SB1_n680) );
  NOR2_X1 R2_SB_SB1_U392 ( .A1(R2_SB_n339), .A2(R2_SB_n341), .ZN(
        R2_SB_SB1_n646) );
  NAND2_X1 R2_SB_SB1_U391 ( .A1(R2_SB_n342), .A2(R2_SB_SB1_n872), .ZN(
        R2_SB_SB1_n770) );
  NOR2_X1 R2_SB_SB1_U390 ( .A1(R2_SB_SB1_n895), .A2(R2_SB_n340), .ZN(
        R2_SB_SB1_n783) );
  NOR2_X1 R2_SB_SB1_U389 ( .A1(R2_SB_n341), .A2(R2_SB_n342), .ZN(
        R2_SB_SB1_n617) );
  NOR2_X1 R2_SB_SB1_U388 ( .A1(R2_SB_SB1_n854), .A2(R2_SB_n339), .ZN(
        R2_SB_SB1_n811) );
  INV_X1 R2_SB_SB1_U387 ( .A(R2_SB_n344), .ZN(R2_SB_SB1_n881) );
  AOI22_X1 R2_SB_SB1_U386 ( .A1(R2_SB_n339), .A2(R2_SB_SB1_n638), .B1(
        R2_SB_SB1_n795), .B2(R2_SB_SB1_n713), .ZN(R2_SB_SB1_n711) );
  NOR2_X1 R2_SB_SB1_U385 ( .A1(R2_SB_SB1_n854), .A2(R2_SB_n342), .ZN(
        R2_SB_SB1_n694) );
  NAND2_X1 R2_SB_SB1_U384 ( .A1(R2_SB_n339), .A2(R2_SB_n342), .ZN(
        R2_SB_SB1_n608) );
  OAI221_X1 R2_SB_SB1_U383 ( .B1(R2_SB_n339), .B2(R2_SB_SB1_n551), .C1(
        R2_SB_SB1_n550), .C2(R2_SB_SB1_n910), .A(R2_SB_SB1_n902), .ZN(
        R2_SB_SB1_n552) );
  OAI221_X1 R2_SB_SB1_U382 ( .B1(R2_SB_SB1_n864), .B2(R2_SB_SB1_n838), .C1(
        R2_SB_SB1_n827), .C2(R2_SB_SB1_n849), .A(R2_SB_SB1_n615), .ZN(
        R2_SB_SB1_n553) );
  OAI221_X1 R2_SB_SB1_U381 ( .B1(R2_SB_SB1_n864), .B2(R2_SB_SB1_n835), .C1(
        R2_SB_SB1_n832), .C2(R2_SB_SB1_n853), .A(R2_SB_SB1_n546), .ZN(
        R2_SB_SB1_n554) );
  AOI221_X1 R2_SB_SB1_U380 ( .B1(R2_SB_SB1_n752), .B2(R2_SB_SB1_n554), .C1(
        R2_SB_SB1_n702), .C2(R2_SB_SB1_n553), .A(R2_SB_SB1_n552), .ZN(
        R2_SB_SB1_n559) );
  OAI22_X1 R2_SB_SB1_U379 ( .A1(R2_SB_SB1_n583), .A2(R2_SB_SB1_n826), .B1(
        R2_SB_SB1_n838), .B2(R2_SB_SB1_n891), .ZN(R2_SB_SB1_n584) );
  OAI211_X1 R2_SB_SB1_U378 ( .C1(R2_SB_SB1_n453), .C2(R2_SB_SB1_n844), .A(
        R2_SB_SB1_n835), .B(R2_SB_SB1_n847), .ZN(R2_SB_SB1_n585) );
  OAI211_X1 R2_SB_SB1_U377 ( .C1(R2_SB_n337), .C2(R2_SB_SB1_n898), .A(
        R2_SB_SB1_n582), .B(R2_SB_SB1_n581), .ZN(R2_SB_SB1_n586) );
  AOI221_X1 R2_SB_SB1_U376 ( .B1(R2_SB_n339), .B2(R2_SB_SB1_n586), .C1(
        R2_SB_SB1_n755), .C2(R2_SB_SB1_n585), .A(R2_SB_SB1_n584), .ZN(
        R2_SB_SB1_n599) );
  OAI221_X1 R2_SB_SB1_U375 ( .B1(R2_SB_SB1_n840), .B2(R2_SB_SB1_n859), .C1(
        R2_SB_SB1_n863), .C2(R2_SB_SB1_n834), .A(R2_SB_SB1_n574), .ZN(
        R2_SB_SB1_n580) );
  OAI22_X1 R2_SB_SB1_U374 ( .A1(R2_SB_n340), .A2(R2_SB_SB1_n578), .B1(
        R2_SB_SB1_n577), .B2(R2_SB_SB1_n831), .ZN(R2_SB_SB1_n579) );
  INV_X1 R2_SB_SB1_U373 ( .A(R2_SB_SB1_n573), .ZN(R2_SB_SB1_n889) );
  AOI221_X1 R2_SB_SB1_U372 ( .B1(R2_SB_SB1_n889), .B2(R2_SB_SB1_n696), .C1(
        R2_SB_SB1_n752), .C2(R2_SB_SB1_n580), .A(R2_SB_SB1_n579), .ZN(
        R2_SB_SB1_n600) );
  NOR2_X1 R2_SB_SB1_U371 ( .A1(R2_SB_n340), .A2(R2_SB_n341), .ZN(
        R2_SB_SB1_n656) );
  INV_X1 R2_SB_SB1_U370 ( .A(R2_SB_n343), .ZN(R2_SB_SB1_n872) );
  NOR3_X1 R2_SB_SB1_U369 ( .A1(R2_SB_SB1_n850), .A2(R2_SB_n341), .A3(
        R2_SB_SB1_n881), .ZN(R2_SB_SB1_n556) );
  NOR2_X1 R2_SB_SB1_U368 ( .A1(R2_SB_SB1_n830), .A2(R2_SB_n341), .ZN(
        R2_SB_SB1_n678) );
  AOI221_X1 R2_SB_SB1_U367 ( .B1(R2_SB_SB1_n806), .B2(R2_SB_SB1_n89), .C1(
        R2_SB_SB1_n805), .C2(R2_SB_SB1_n804), .A(R2_SB_SB1_n803), .ZN(
        R2_SB_SB1_n807) );
  AOI211_X1 R2_SB_SB1_U366 ( .C1(R2_SB_SB1_n799), .C2(R2_SB_SB1_n798), .A(
        R2_SB_SB1_n797), .B(R2_SB_SB1_n796), .ZN(R2_SB_SB1_n808) );
  AOI22_X1 R2_SB_SB1_U365 ( .A1(R2_SB_SB1_n793), .A2(R2_SB_SB1_n792), .B1(
        R2_SB_SB1_n791), .B2(R2_SB_SB1_n790), .ZN(R2_SB_SB1_n809) );
  OAI221_X1 R2_SB_SB1_U364 ( .B1(R2_SB_n343), .B2(R2_SB_SB1_n809), .C1(
        R2_SB_SB1_n808), .C2(R2_SB_SB1_n859), .A(R2_SB_SB1_n807), .ZN(
        R2_SB_SB1_n821) );
  NOR2_X1 R2_SB_SB1_U363 ( .A1(R2_SB_n344), .A2(R2_SB_n341), .ZN(
        R2_SB_SB1_n489) );
  OAI21_X1 R2_SB_SB1_U362 ( .B1(R2_SB_SB1_n864), .B2(R2_SB_SB1_n878), .A(
        R2_SB_SB1_n894), .ZN(R2_SB_SB1_n490) );
  AOI221_X1 R2_SB_SB1_U361 ( .B1(R2_SB_SB1_n779), .B2(R2_SB_SB1_n490), .C1(
        R2_SB_SB1_n489), .C2(R2_SB_SB1_n782), .A(R2_SB_SB1_n756), .ZN(
        R2_SB_SB1_n491) );
  AOI222_X1 R2_SB_SB1_U360 ( .A1(R2_SB_SB1_n789), .A2(R2_SB_SB1_n772), .B1(
        R2_SB_SB1_n646), .B2(R2_SB_SB1_n813), .C1(R2_SB_SB1_n709), .C2(
        R2_SB_SB1_n811), .ZN(R2_SB_SB1_n647) );
  OAI221_X1 R2_SB_SB1_U359 ( .B1(R2_SB_n338), .B2(R2_SB_SB1_n884), .C1(
        R2_SB_SB1_n453), .C2(R2_SB_SB1_n880), .A(R2_SB_SB1_n649), .ZN(
        R2_SB_SB1_n650) );
  OAI221_X1 R2_SB_SB1_U358 ( .B1(R2_SB_n340), .B2(R2_SB_SB1_n648), .C1(
        R2_SB_SB1_n845), .C2(R2_SB_SB1_n868), .A(R2_SB_SB1_n647), .ZN(
        R2_SB_SB1_n652) );
  AOI222_X1 R2_SB_SB1_U357 ( .A1(R2_SB_SB1_n781), .A2(R2_SB_SB1_n652), .B1(
        R2_SB_SB1_n651), .B2(R2_SB_SB1_n730), .C1(R2_SB_SB1_n782), .C2(
        R2_SB_SB1_n650), .ZN(R2_SB_SB1_n693) );
  NOR2_X1 R2_SB_SB1_U356 ( .A1(R2_SB_SB1_n863), .A2(R2_SB_n340), .ZN(
        R2_SB_SB1_n618) );
  NOR3_X1 R2_SB_SB1_U355 ( .A1(R2_SB_SB1_n840), .A2(R2_SB_n343), .A3(
        R2_SB_SB1_n869), .ZN(R2_SB_SB1_n575) );
  AOI221_X1 R2_SB_SB1_U354 ( .B1(R2_SB_SB1_n591), .B2(R2_SB_SB1_n453), .C1(
        R2_SB_SB1_n576), .C2(R2_SB_SB1_n684), .A(R2_SB_SB1_n575), .ZN(
        R2_SB_SB1_n578) );
  OAI211_X1 R2_SB_SB1_U353 ( .C1(R2_SB_n342), .C2(R2_SB_SB1_n848), .A(
        R2_SB_SB1_n860), .B(R2_SB_SB1_n853), .ZN(R2_SB_SB1_n662) );
  OAI21_X1 R2_SB_SB1_U352 ( .B1(R2_SB_SB1_n876), .B2(R2_SB_SB1_n853), .A(
        R2_SB_SB1_n908), .ZN(R2_SB_SB1_n663) );
  AOI221_X1 R2_SB_SB1_U351 ( .B1(R2_SB_SB1_n779), .B2(R2_SB_SB1_n663), .C1(
        R2_SB_SB1_n702), .C2(R2_SB_SB1_n662), .A(R2_SB_SB1_n661), .ZN(
        R2_SB_SB1_n664) );
  OAI222_X1 R2_SB_SB1_U350 ( .A1(R2_SB_SB1_n718), .A2(R2_SB_SB1_n907), .B1(
        R2_SB_SB1_n452), .B2(R2_SB_SB1_n664), .C1(R2_SB_SB1_n832), .C2(
        R2_SB_SB1_n802), .ZN(R2_SB_SB1_n667) );
  NOR3_X1 R2_SB_SB1_U349 ( .A1(R2_SB_SB1_n849), .A2(R2_SB_n344), .A3(
        R2_SB_SB1_n854), .ZN(R2_SB_SB1_n605) );
  OAI22_X1 R2_SB_SB1_U348 ( .A1(R2_SB_n343), .A2(R2_SB_n341), .B1(R2_SB_n342), 
        .B2(R2_SB_SB1_n883), .ZN(R2_SB_SB1_n606) );
  AOI221_X1 R2_SB_SB1_U347 ( .B1(R2_SB_SB1_n755), .B2(R2_SB_SB1_n791), .C1(
        R2_SB_SB1_n758), .C2(R2_SB_SB1_n606), .A(R2_SB_SB1_n605), .ZN(
        R2_SB_SB1_n607) );
  NOR2_X1 R2_SB_SB1_U346 ( .A1(R2_SB_SB1_n452), .A2(R2_SB_n339), .ZN(
        R2_SB_SB1_n794) );
  NOR2_X1 R2_SB_SB1_U345 ( .A1(R2_SB_n342), .A2(R2_SB_n344), .ZN(
        R2_SB_SB1_n709) );
  NOR2_X1 R2_SB_SB1_U344 ( .A1(R2_SB_SB1_n830), .A2(R2_SB_n340), .ZN(
        R2_SB_SB1_n782) );
  NOR3_X1 R2_SB_SB1_U343 ( .A1(R2_SB_SB1_n901), .A2(R2_SB_n343), .A3(
        R2_SB_SB1_n843), .ZN(R2_SB_SB1_n729) );
  AOI221_X1 R2_SB_SB1_U342 ( .B1(R2_SB_SB1_n805), .B2(R2_SB_SB1_n813), .C1(
        R2_SB_SB1_n789), .C2(R2_SB_SB1_n728), .A(R2_SB_SB1_n727), .ZN(
        R2_SB_SB1_n732) );
  AOI211_X1 R2_SB_SB1_U341 ( .C1(R2_SB_SB1_n752), .C2(R2_SB_SB1_n730), .A(
        R2_SB_SB1_n759), .B(R2_SB_SB1_n729), .ZN(R2_SB_SB1_n731) );
  OAI222_X1 R2_SB_SB1_U340 ( .A1(R2_SB_SB1_n733), .A2(R2_SB_SB1_n839), .B1(
        R2_SB_SB1_n732), .B2(R2_SB_SB1_n837), .C1(R2_SB_SB1_n731), .C2(
        R2_SB_SB1_n835), .ZN(R2_SB_SB1_n734) );
  NOR2_X1 R2_SB_SB1_U339 ( .A1(R2_SB_SB1_n854), .A2(R2_SB_n340), .ZN(
        R2_SB_SB1_n805) );
  NOR2_X1 R2_SB_SB1_U338 ( .A1(R2_SB_SB1_n872), .A2(R2_SB_n342), .ZN(
        R2_SB_SB1_n767) );
  INV_X1 R2_SB_SB1_U337 ( .A(R2_SB_n339), .ZN(R2_SB_SB1_n830) );
  NOR2_X1 R2_SB_SB1_U336 ( .A1(R2_SB_n343), .A2(R2_SB_n344), .ZN(
        R2_SB_SB1_n702) );
  NOR2_X1 R2_SB_SB1_U335 ( .A1(R2_SB_n338), .A2(R2_SB_n339), .ZN(
        R2_SB_SB1_n795) );
  NOR2_X1 R2_SB_SB1_U334 ( .A1(R2_SB_n342), .A2(R2_SB_n343), .ZN(
        R2_SB_SB1_n813) );
  NOR3_X1 R2_SB_SB1_U333 ( .A1(R2_SB_SB1_n833), .A2(R2_SB_n340), .A3(
        R2_SB_SB1_n885), .ZN(R2_SB_SB1_n639) );
  INV_X1 R2_SB_SB1_U332 ( .A(R2_SB_n341), .ZN(R2_SB_SB1_n854) );
  NOR2_X1 R2_SB_SB1_U331 ( .A1(R2_SB_SB1_n843), .A2(R2_SB_n339), .ZN(
        R2_SB_SB1_n792) );
  INV_X1 R2_SB_SB1_U330 ( .A(R2_SB_n342), .ZN(R2_SB_SB1_n863) );
  NAND2_X1 R2_SB_SB1_U329 ( .A1(R2_SB_SB1_n791), .A2(R2_SB_SB1_n772), .ZN(
        R2_SB_SB1_n775) );
  OAI21_X1 R2_SB_SB1_U328 ( .B1(R2_SB_SB1_n775), .B2(R2_SB_SB1_n774), .A(
        R2_SB_SB1_n773), .ZN(R2_SB_SB1_n776) );
  INV_X1 R2_SB_SB1_U327 ( .A(R2_SB_SB1_n776), .ZN(R2_SB_SB1_n887) );
  INV_X1 R2_SB_SB1_U326 ( .A(R2_SB_SB1_n783), .ZN(R2_SB_SB1_n897) );
  INV_X1 R2_SB_SB1_U325 ( .A(R2_SB_SB1_n678), .ZN(R2_SB_SB1_n860) );
  INV_X1 R2_SB_SB1_U324 ( .A(R2_SB_SB1_n811), .ZN(R2_SB_SB1_n855) );
  INV_X1 R2_SB_SB1_U323 ( .A(R2_SB_SB1_n463), .ZN(R2_SB_SB1_n842) );
  INV_X1 R2_SB_SB1_U322 ( .A(R2_SB_SB1_n711), .ZN(R2_SB_SB1_n909) );
  NAND2_X1 R2_SB_SB1_U321 ( .A1(R2_SB_SB1_n678), .A2(R2_SB_SB1_n781), .ZN(
        R2_SB_SB1_n615) );
  NAND2_X1 R2_SB_SB1_U320 ( .A1(R2_SB_SB1_n680), .A2(R2_SB_SB1_n810), .ZN(
        R2_SB_SB1_n581) );
  NAND2_X1 R2_SB_SB1_U319 ( .A1(R2_SB_SB1_n772), .A2(R2_SB_SB1_n684), .ZN(
        R2_SB_SB1_n785) );
  NAND2_X1 R2_SB_SB1_U318 ( .A1(R2_SB_SB1_n670), .A2(R2_SB_SB1_n881), .ZN(
        R2_SB_SB1_n773) );
  NAND2_X1 R2_SB_SB1_U317 ( .A1(R2_SB_SB1_n670), .A2(R2_SB_SB1_n872), .ZN(
        R2_SB_SB1_n801) );
  NAND2_X1 R2_SB_SB1_U316 ( .A1(R2_SB_SB1_n452), .A2(R2_SB_SB1_n843), .ZN(
        R2_SB_SB1_n548) );
  NOR2_X1 R2_SB_SB1_U315 ( .A1(R2_SB_SB1_n854), .A2(R2_SB_SB1_n827), .ZN(
        R2_SB_SB1_n793) );
  OAI21_X1 R2_SB_SB1_U314 ( .B1(R2_SB_SB1_n718), .B2(R2_SB_SB1_n588), .A(
        R2_SB_SB1_n587), .ZN(R2_SB_SB1_n597) );
  AOI22_X1 R2_SB_SB1_U313 ( .A1(R2_SB_SB1_n753), .A2(R2_SB_SB1_n771), .B1(
        R2_SB_SB1_n752), .B2(R2_SB_SB1_n751), .ZN(R2_SB_SB1_n825) );
  AOI22_X1 R2_SB_SB1_U312 ( .A1(R2_SB_n338), .A2(R2_SB_SB1_n765), .B1(
        R2_SB_SB1_n764), .B2(R2_SB_SB1_n453), .ZN(R2_SB_SB1_n824) );
  NOR4_X1 R2_SB_SB1_U311 ( .A1(R2_SB_SB1_n464), .A2(R2_SB_SB1_n886), .A3(
        R2_SB_SB1_n555), .A4(R2_SB_SB1_n639), .ZN(R2_SB_SB1_n486) );
  AOI211_X1 R2_SB_SB1_U310 ( .C1(R2_SB_SB1_n684), .C2(R2_SB_SB1_n462), .A(
        R2_SB_SB1_n461), .B(R2_SB_SB1_n460), .ZN(R2_SB_SB1_n487) );
  AOI221_X1 R2_SB_SB1_U309 ( .B1(R2_SB_SB1_n810), .B2(R2_SB_SB1_n533), .C1(
        R2_SB_SB1_n565), .C2(R2_SB_n338), .A(R2_SB_SB1_n532), .ZN(
        R2_SB_SB1_n561) );
  NOR4_X1 R2_SB_SB1_U308 ( .A1(R2_SB_SB1_n557), .A2(R2_SB_SB1_n556), .A3(
        R2_SB_SB1_n555), .A4(R2_SB_SB1_n674), .ZN(R2_SB_SB1_n558) );
  AOI221_X1 R2_SB_SB1_U307 ( .B1(R2_SB_SB1_n772), .B2(R2_SB_SB1_n572), .C1(
        R2_SB_SB1_n753), .C2(R2_SB_SB1_n758), .A(R2_SB_SB1_n571), .ZN(
        R2_SB_SB1_n601) );
  AOI211_X1 R2_SB_SB1_U306 ( .C1(R2_SB_SB1_n597), .C2(R2_SB_SB1_n453), .A(
        R2_SB_SB1_n596), .B(R2_SB_SB1_n595), .ZN(R2_SB_SB1_n598) );
  AOI221_X1 R2_SB_SB1_U305 ( .B1(R2_SB_SB1_n604), .B2(R2_SB_SB1_n877), .C1(
        R2_SB_SB1_n603), .C2(R2_SB_SB1_n679), .A(R2_SB_SB1_n602), .ZN(
        R2_SB_SB1_n645) );
  NOR4_X1 R2_SB_SB1_U304 ( .A1(R2_SB_SB1_n641), .A2(R2_SB_SB1_n640), .A3(
        R2_SB_SB1_n639), .A4(R2_SB_SB1_n673), .ZN(R2_SB_SB1_n642) );
  OAI21_X1 R2_SB_SB1_U303 ( .B1(R2_SB_SB1_n810), .B2(R2_SB_SB1_n744), .A(
        R2_SB_SB1_n743), .ZN(R2_SB_SB1_n745) );
  NOR4_X1 R2_SB_SB1_U302 ( .A1(R2_SB_SB1_n737), .A2(R2_SB_SB1_n736), .A3(
        R2_SB_SB1_n735), .A4(R2_SB_SB1_n734), .ZN(R2_SB_SB1_n738) );
  AOI211_X1 R2_SB_SB1_U301 ( .C1(R2_SB_SB1_n713), .C2(R2_SB_SB1_n758), .A(
        R2_SB_SB1_n712), .B(R2_SB_SB1_n909), .ZN(R2_SB_SB1_n739) );
  NOR4_X1 R2_SB_SB1_U300 ( .A1(R2_SB_SB1_n689), .A2(R2_SB_SB1_n688), .A3(
        R2_SB_SB1_n687), .A4(R2_SB_SB1_n686), .ZN(R2_SB_SB1_n690) );
  AOI211_X1 R2_SB_SB1_U299 ( .C1(R2_SB_SB1_n752), .C2(R2_SB_SB1_n668), .A(
        R2_SB_SB1_n667), .B(R2_SB_SB1_n666), .ZN(R2_SB_SB1_n691) );
  AOI221_X1 R2_SB_SB1_U298 ( .B1(R2_SB_SB1_n565), .B2(R2_SB_SB1_n766), .C1(
        R2_SB_SB1_n759), .C2(R2_SB_SB1_n791), .A(R2_SB_SB1_n513), .ZN(
        R2_SB_SB1_n525) );
  NOR4_X1 R2_SB_SB1_U297 ( .A1(R2_SB_SB1_n523), .A2(R2_SB_SB1_n522), .A3(
        R2_SB_SB1_n521), .A4(R2_SB_SB1_n520), .ZN(R2_SB_SB1_n524) );
  OAI221_X1 R2_SB_SB1_U296 ( .B1(R2_SB_SB1_n849), .B2(R2_SB_SB1_n770), .C1(
        R2_SB_SB1_n883), .C2(R2_SB_SB1_n608), .A(R2_SB_SB1_n567), .ZN(
        R2_SB_SB1_n568) );
  OAI21_X1 R2_SB_SB1_U295 ( .B1(R2_SB_SB1_n569), .B2(R2_SB_SB1_n568), .A(
        R2_SB_SB1_n781), .ZN(R2_SB_SB1_n570) );
  OAI21_X1 R2_SB_SB1_U294 ( .B1(R2_SB_SB1_n839), .B2(R2_SB_SB1_n892), .A(
        R2_SB_SB1_n570), .ZN(R2_SB_SB1_n571) );
  INV_X1 R2_SB_SB1_U293 ( .A(R2_SB_SB1_n780), .ZN(R2_SB_SB1_n870) );
  OAI21_X1 R2_SB_SB1_U292 ( .B1(R2_SB_SB1_n778), .B2(R2_SB_SB1_n744), .A(
        R2_SB_SB1_n696), .ZN(R2_SB_SB1_n508) );
  OAI211_X1 R2_SB_SB1_U291 ( .C1(R2_SB_SB1_n813), .C2(R2_SB_SB1_n812), .A(
        R2_SB_SB1_n811), .B(R2_SB_SB1_n810), .ZN(R2_SB_SB1_n817) );
  INV_X1 R2_SB_SB1_U290 ( .A(R2_SB_SB1_n743), .ZN(R2_SB_SB1_n851) );
  AND3_X1 R2_SB_SB1_U289 ( .A1(R2_SB_SB1_n779), .A2(R2_SB_SB1_n812), .A3(
        R2_SB_SB1_n656), .ZN(R2_SB_SB1_n87) );
  NOR3_X1 R2_SB_SB1_U288 ( .A1(R2_SB_SB1_n858), .A2(R2_SB_SB1_n665), .A3(
        R2_SB_SB1_n890), .ZN(R2_SB_SB1_n13) );
  OR3_X1 R2_SB_SB1_U287 ( .A1(R2_SB_SB1_n13), .A2(R2_SB_SB1_n675), .A3(
        R2_SB_SB1_n87), .ZN(R2_SB_SB1_n464) );
  OAI22_X1 R2_SB_SB1_U286 ( .A1(R2_SB_SB1_n872), .A2(R2_SB_SB1_n857), .B1(
        R2_SB_SB1_n854), .B2(R2_SB_SB1_n876), .ZN(R2_SB_SB1_n547) );
  INV_X1 R2_SB_SB1_U285 ( .A(R2_SB_SB1_n582), .ZN(R2_SB_SB1_n911) );
  AOI21_X1 R2_SB_SB1_U284 ( .B1(R2_SB_SB1_n781), .B2(R2_SB_SB1_n547), .A(
        R2_SB_SB1_n911), .ZN(R2_SB_SB1_n551) );
  AOI21_X1 R2_SB_SB1_U283 ( .B1(R2_SB_SB1_n754), .B2(R2_SB_SB1_n758), .A(
        R2_SB_SB1_n467), .ZN(R2_SB_SB1_n468) );
  AOI21_X1 R2_SB_SB1_U282 ( .B1(R2_SB_SB1_n778), .B2(R2_SB_SB1_n453), .A(
        R2_SB_SB1_n789), .ZN(R2_SB_SB1_n700) );
  AOI22_X1 R2_SB_SB1_U281 ( .A1(R2_SB_SB1_n725), .A2(R2_SB_SB1_n617), .B1(
        R2_SB_SB1_n766), .B2(R2_SB_SB1_n730), .ZN(R2_SB_SB1_n562) );
  AOI21_X1 R2_SB_SB1_U280 ( .B1(R2_SB_SB1_n743), .B2(R2_SB_n338), .A(
        R2_SB_SB1_n747), .ZN(R2_SB_SB1_n564) );
  OAI21_X1 R2_SB_SB1_U279 ( .B1(R2_SB_SB1_n684), .B2(R2_SB_SB1_n799), .A(
        R2_SB_SB1_n780), .ZN(R2_SB_SB1_n563) );
  OAI211_X1 R2_SB_SB1_U278 ( .C1(R2_SB_SB1_n564), .C2(R2_SB_SB1_n868), .A(
        R2_SB_SB1_n563), .B(R2_SB_SB1_n562), .ZN(R2_SB_SB1_n572) );
  OAI21_X1 R2_SB_SB1_U277 ( .B1(R2_SB_SB1_n905), .B2(R2_SB_SB1_n859), .A(
        R2_SB_SB1_n895), .ZN(R2_SB_SB1_n529) );
  AOI211_X1 R2_SB_SB1_U276 ( .C1(R2_SB_SB1_n529), .C2(R2_SB_SB1_n830), .A(
        R2_SB_SB1_n633), .B(R2_SB_SB1_n528), .ZN(R2_SB_SB1_n530) );
  AOI22_X1 R2_SB_SB1_U275 ( .A1(R2_SB_SB1_n680), .A2(R2_SB_SB1_n843), .B1(
        R2_SB_SB1_n678), .B2(R2_SB_SB1_n772), .ZN(R2_SB_SB1_n531) );
  OAI211_X1 R2_SB_SB1_U274 ( .C1(R2_SB_SB1_n905), .C2(R2_SB_SB1_n864), .A(
        R2_SB_SB1_n531), .B(R2_SB_SB1_n530), .ZN(R2_SB_SB1_n533) );
  OAI21_X1 R2_SB_SB1_U273 ( .B1(R2_SB_SB1_n755), .B2(R2_SB_SB1_n754), .A(
        R2_SB_SB1_n782), .ZN(R2_SB_SB1_n757) );
  INV_X1 R2_SB_SB1_U272 ( .A(R2_SB_SB1_n756), .ZN(R2_SB_SB1_n899) );
  OAI211_X1 R2_SB_SB1_U271 ( .C1(R2_SB_SB1_n845), .C2(R2_SB_SB1_n880), .A(
        R2_SB_SB1_n757), .B(R2_SB_SB1_n899), .ZN(R2_SB_SB1_n765) );
  INV_X1 R2_SB_SB1_U270 ( .A(R2_SB_SB1_n696), .ZN(R2_SB_SB1_n836) );
  AOI21_X1 R2_SB_SB1_U269 ( .B1(R2_SB_SB1_n843), .B2(R2_SB_SB1_n835), .A(
        R2_SB_SB1_n879), .ZN(R2_SB_SB1_n595) );
  NAND2_X1 R2_SB_SB1_U268 ( .A1(R2_SB_SB1_n634), .A2(R2_SB_SB1_n805), .ZN(
        R2_SB_SB1_n800) );
  NAND2_X1 R2_SB_SB1_U267 ( .A1(R2_SB_SB1_n772), .A2(R2_SB_SB1_n507), .ZN(
        R2_SB_SB1_n648) );
  AOI21_X1 R2_SB_SB1_U266 ( .B1(R2_SB_SB1_n849), .B2(R2_SB_SB1_n608), .A(
        R2_SB_SB1_n878), .ZN(R2_SB_SB1_n528) );
  INV_X1 R2_SB_SB1_U265 ( .A(R2_SB_SB1_n794), .ZN(R2_SB_SB1_n837) );
  NOR2_X1 R2_SB_SB1_U263 ( .A1(R2_SB_SB1_n770), .A2(R2_SB_SB1_n833), .ZN(
        R2_SB_SB1_n651) );
  INV_X1 R2_SB_SB1_U262 ( .A(R2_SB_SB1_n798), .ZN(R2_SB_SB1_n901) );
  INV_X1 R2_SB_SB1_U261 ( .A(R2_SB_SB1_n813), .ZN(R2_SB_SB1_n876) );
  AOI22_X1 R2_SB_SB1_U260 ( .A1(R2_SB_SB1_n696), .A2(R2_SB_SB1_n789), .B1(
        R2_SB_SB1_n778), .B2(R2_SB_SB1_n779), .ZN(R2_SB_SB1_n612) );
  AOI22_X1 R2_SB_SB1_U259 ( .A1(R2_SB_SB1_n795), .A2(R2_SB_SB1_n798), .B1(
        R2_SB_SB1_n767), .B2(R2_SB_SB1_n766), .ZN(R2_SB_SB1_n768) );
  NAND2_X1 R2_SB_SB1_U258 ( .A1(R2_SB_SB1_n865), .A2(R2_SB_SB1_n853), .ZN(
        R2_SB_SB1_n495) );
  AOI22_X1 R2_SB_SB1_U257 ( .A1(R2_SB_SB1_n684), .A2(R2_SB_SB1_n495), .B1(
        R2_SB_SB1_n696), .B2(R2_SB_SB1_n618), .ZN(R2_SB_SB1_n496) );
  INV_X1 R2_SB_SB1_U256 ( .A(R2_SB_SB1_n805), .ZN(R2_SB_SB1_n857) );
  NAND2_X1 R2_SB_SB1_U255 ( .A1(R2_SB_SB1_n843), .A2(R2_SB_SB1_n863), .ZN(
        R2_SB_SB1_n774) );
  AOI22_X1 R2_SB_SB1_U254 ( .A1(R2_SB_SB1_n798), .A2(R2_SB_SB1_n627), .B1(
        R2_SB_SB1_n743), .B2(R2_SB_SB1_n752), .ZN(R2_SB_SB1_n567) );
  INV_X1 R2_SB_SB1_U253 ( .A(R2_SB_SB1_n767), .ZN(R2_SB_SB1_n874) );
  NOR2_X1 R2_SB_SB1_U252 ( .A1(R2_SB_SB1_n795), .A2(R2_SB_SB1_n794), .ZN(
        R2_SB_SB1_n814) );
  INV_X1 R2_SB_SB1_U251 ( .A(R2_SB_SB1_n694), .ZN(R2_SB_SB1_n869) );
  NOR2_X1 R2_SB_SB1_U250 ( .A1(R2_SB_SB1_n830), .A2(R2_SB_SB1_n684), .ZN(
        R2_SB_SB1_n665) );
  NOR2_X1 R2_SB_SB1_U249 ( .A1(R2_SB_SB1_n843), .A2(R2_SB_n338), .ZN(
        R2_SB_SB1_n604) );
  NOR2_X1 R2_SB_SB1_U248 ( .A1(R2_SB_SB1_n863), .A2(R2_SB_SB1_n858), .ZN(
        R2_SB_SB1_n790) );
  NAND2_X1 R2_SB_SB1_U247 ( .A1(R2_SB_SB1_n752), .A2(R2_SB_SB1_n507), .ZN(
        R2_SB_SB1_n802) );
  AOI21_X1 R2_SB_SB1_U246 ( .B1(R2_SB_SB1_n789), .B2(R2_SB_SB1_n798), .A(
        R2_SB_SB1_n783), .ZN(R2_SB_SB1_n721) );
  OAI21_X1 R2_SB_SB1_U245 ( .B1(R2_SB_SB1_n747), .B2(R2_SB_SB1_n843), .A(
        R2_SB_SB1_n759), .ZN(R2_SB_SB1_n719) );
  OR3_X1 R2_SB_SB1_U244 ( .A1(R2_SB_SB1_n718), .A2(R2_SB_SB1_n452), .A3(
        R2_SB_SB1_n802), .ZN(R2_SB_SB1_n720) );
  OAI211_X1 R2_SB_SB1_U243 ( .C1(R2_SB_SB1_n721), .C2(R2_SB_SB1_n826), .A(
        R2_SB_SB1_n720), .B(R2_SB_SB1_n719), .ZN(R2_SB_SB1_n736) );
  AOI22_X1 R2_SB_SB1_U242 ( .A1(R2_SB_SB1_n678), .A2(R2_SB_SB1_n767), .B1(
        R2_SB_SB1_n900), .B2(R2_SB_SB1_n843), .ZN(R2_SB_SB1_n683) );
  OAI21_X1 R2_SB_SB1_U241 ( .B1(R2_SB_SB1_n794), .B2(R2_SB_SB1_n791), .A(
        R2_SB_SB1_n882), .ZN(R2_SB_SB1_n681) );
  OAI21_X1 R2_SB_SB1_U240 ( .B1(R2_SB_SB1_n680), .B2(R2_SB_SB1_n679), .A(
        R2_SB_SB1_n696), .ZN(R2_SB_SB1_n682) );
  OAI211_X1 R2_SB_SB1_U239 ( .C1(R2_SB_SB1_n683), .C2(R2_SB_SB1_n829), .A(
        R2_SB_SB1_n682), .B(R2_SB_SB1_n681), .ZN(R2_SB_SB1_n688) );
  NOR3_X1 R2_SB_SB1_U238 ( .A1(R2_SB_SB1_n848), .A2(R2_SB_SB1_n452), .A3(
        R2_SB_SB1_n863), .ZN(R2_SB_SB1_n540) );
  OAI22_X1 R2_SB_SB1_U237 ( .A1(R2_SB_SB1_n858), .A2(R2_SB_SB1_n838), .B1(
        R2_SB_SB1_n857), .B2(R2_SB_SB1_n840), .ZN(R2_SB_SB1_n541) );
  AOI21_X1 R2_SB_SB1_U236 ( .B1(R2_SB_n338), .B2(R2_SB_SB1_n548), .A(
        R2_SB_SB1_n862), .ZN(R2_SB_SB1_n539) );
  NOR3_X1 R2_SB_SB1_U235 ( .A1(R2_SB_SB1_n541), .A2(R2_SB_SB1_n540), .A3(
        R2_SB_SB1_n539), .ZN(R2_SB_SB1_n542) );
  AOI21_X1 R2_SB_SB1_U234 ( .B1(R2_SB_SB1_n730), .B2(R2_SB_SB1_n709), .A(
        R2_SB_SB1_n753), .ZN(R2_SB_SB1_n733) );
  INV_X1 R2_SB_SB1_U233 ( .A(R2_SB_SB1_n791), .ZN(R2_SB_SB1_n840) );
  NOR3_X1 R2_SB_SB1_U232 ( .A1(R2_SB_SB1_n828), .A2(R2_SB_SB1_n856), .A3(
        R2_SB_SB1_n876), .ZN(R2_SB_SB1_n819) );
  AOI21_X1 R2_SB_SB1_U231 ( .B1(R2_SB_SB1_n845), .B2(R2_SB_SB1_n837), .A(
        R2_SB_SB1_n906), .ZN(R2_SB_SB1_n818) );
  NOR4_X1 R2_SB_SB1_U230 ( .A1(R2_SB_SB1_n821), .A2(R2_SB_SB1_n820), .A3(
        R2_SB_SB1_n819), .A4(R2_SB_SB1_n818), .ZN(R2_SB_SB1_n822) );
  INV_X1 R2_SB_SB1_U229 ( .A(R2_SB_SB1_n789), .ZN(R2_SB_SB1_n853) );
  NOR2_X1 R2_SB_SB1_U228 ( .A1(R2_SB_SB1_n743), .A2(R2_SB_SB1_n603), .ZN(
        R2_SB_SB1_n718) );
  AOI221_X1 R2_SB_SB1_U227 ( .B1(R2_SB_SB1_n877), .B2(R2_SB_SB1_n684), .C1(
        R2_SB_SB1_n591), .C2(R2_SB_SB1_n89), .A(R2_SB_SB1_n590), .ZN(
        R2_SB_SB1_n593) );
  AOI22_X1 R2_SB_SB1_U226 ( .A1(R2_SB_SB1_n810), .A2(R2_SB_SB1_n589), .B1(
        R2_SB_SB1_n798), .B2(R2_SB_SB1_n723), .ZN(R2_SB_SB1_n594) );
  OAI221_X1 R2_SB_SB1_U225 ( .B1(R2_SB_SB1_n594), .B2(R2_SB_SB1_n859), .C1(
        R2_SB_SB1_n593), .C2(R2_SB_SB1_n849), .A(R2_SB_SB1_n592), .ZN(
        R2_SB_SB1_n596) );
  INV_X1 R2_SB_SB1_U224 ( .A(R2_SB_SB1_n744), .ZN(R2_SB_SB1_n868) );
  OAI21_X1 R2_SB_SB1_U223 ( .B1(R2_SB_SB1_n779), .B2(R2_SB_SB1_n453), .A(
        R2_SB_SB1_n656), .ZN(R2_SB_SB1_n503) );
  NOR2_X1 R2_SB_SB1_U222 ( .A1(R2_SB_SB1_n618), .A2(R2_SB_SB1_n780), .ZN(
        R2_SB_SB1_n504) );
  OAI221_X1 R2_SB_SB1_U221 ( .B1(R2_SB_SB1_n504), .B2(R2_SB_SB1_n840), .C1(
        R2_SB_SB1_n869), .C2(R2_SB_SB1_n852), .A(R2_SB_SB1_n503), .ZN(
        R2_SB_SB1_n505) );
  INV_X1 R2_SB_SB1_U220 ( .A(R2_SB_SB1_n617), .ZN(R2_SB_SB1_n862) );
  AOI21_X1 R2_SB_SB1_U219 ( .B1(R2_SB_SB1_n828), .B2(R2_SB_SB1_n850), .A(
        R2_SB_SB1_n879), .ZN(R2_SB_SB1_n459) );
  AOI221_X1 R2_SB_SB1_U218 ( .B1(R2_SB_SB1_n463), .B2(R2_SB_SB1_n591), .C1(
        R2_SB_SB1_n514), .C2(R2_SB_SB1_n766), .A(R2_SB_SB1_n459), .ZN(
        R2_SB_SB1_n488) );
  OAI222_X1 R2_SB_SB1_U217 ( .A1(R2_SB_SB1_n623), .A2(R2_SB_SB1_n851), .B1(
        R2_SB_SB1_n622), .B2(R2_SB_SB1_n883), .C1(R2_SB_SB1_n621), .C2(
        R2_SB_SB1_n905), .ZN(R2_SB_SB1_n624) );
  OAI221_X1 R2_SB_SB1_U216 ( .B1(R2_SB_SB1_n903), .B2(R2_SB_SB1_n844), .C1(
        R2_SB_SB1_n848), .C2(R2_SB_SB1_n910), .A(R2_SB_SB1_n607), .ZN(
        R2_SB_SB1_n626) );
  OAI211_X1 R2_SB_SB1_U215 ( .C1(R2_SB_SB1_n857), .C2(R2_SB_SB1_n831), .A(
        R2_SB_SB1_n612), .B(R2_SB_SB1_n611), .ZN(R2_SB_SB1_n625) );
  AOI221_X1 R2_SB_SB1_U214 ( .B1(R2_SB_SB1_n452), .B2(R2_SB_SB1_n626), .C1(
        R2_SB_SB1_n752), .C2(R2_SB_SB1_n625), .A(R2_SB_SB1_n624), .ZN(
        R2_SB_SB1_n644) );
  OAI22_X1 R2_SB_SB1_U213 ( .A1(R2_SB_SB1_n733), .A2(R2_SB_SB1_n837), .B1(
        R2_SB_SB1_n842), .B2(R2_SB_SB1_n884), .ZN(R2_SB_SB1_n653) );
  OAI22_X1 R2_SB_SB1_U212 ( .A1(R2_SB_SB1_n858), .A2(R2_SB_SB1_n834), .B1(
        R2_SB_n338), .B2(R2_SB_SB1_n859), .ZN(R2_SB_SB1_n654) );
  OAI21_X1 R2_SB_SB1_U211 ( .B1(R2_SB_SB1_n903), .B2(R2_SB_SB1_n859), .A(
        R2_SB_SB1_n895), .ZN(R2_SB_SB1_n655) );
  AOI221_X1 R2_SB_SB1_U210 ( .B1(R2_SB_SB1_n795), .B2(R2_SB_SB1_n655), .C1(
        R2_SB_SB1_n702), .C2(R2_SB_SB1_n654), .A(R2_SB_SB1_n653), .ZN(
        R2_SB_SB1_n692) );
  AOI221_X1 R2_SB_SB1_U209 ( .B1(R2_SB_SB1_n684), .B2(R2_SB_SB1_n536), .C1(
        R2_SB_SB1_n535), .C2(R2_SB_SB1_n628), .A(R2_SB_SB1_n534), .ZN(
        R2_SB_SB1_n537) );
  OAI222_X1 R2_SB_SB1_U208 ( .A1(R2_SB_SB1_n543), .A2(R2_SB_SB1_n847), .B1(
        R2_SB_SB1_n835), .B2(R2_SB_SB1_n573), .C1(R2_SB_SB1_n542), .C2(
        R2_SB_SB1_n883), .ZN(R2_SB_SB1_n544) );
  OAI221_X1 R2_SB_SB1_U207 ( .B1(R2_SB_SB1_n89), .B2(R2_SB_SB1_n588), .C1(
        R2_SB_n337), .C2(R2_SB_SB1_n910), .A(R2_SB_SB1_n537), .ZN(
        R2_SB_SB1_n545) );
  AOI221_X1 R2_SB_SB1_U206 ( .B1(R2_SB_SB1_n792), .B2(R2_SB_SB1_n545), .C1(
        R2_SB_SB1_n753), .C2(R2_SB_SB1_n791), .A(R2_SB_SB1_n544), .ZN(
        R2_SB_SB1_n560) );
  AOI22_X1 R2_SB_SB1_U205 ( .A1(R2_SB_SB1_n798), .A2(R2_SB_SB1_n708), .B1(
        R2_SB_SB1_n795), .B2(R2_SB_SB1_n767), .ZN(R2_SB_SB1_n631) );
  AOI21_X1 R2_SB_SB1_U204 ( .B1(R2_SB_SB1_n755), .B2(R2_SB_SB1_n758), .A(
        R2_SB_SB1_n756), .ZN(R2_SB_SB1_n629) );
  OAI222_X1 R2_SB_SB1_U203 ( .A1(R2_SB_SB1_n631), .A2(R2_SB_SB1_n857), .B1(
        R2_SB_SB1_n630), .B2(R2_SB_SB1_n875), .C1(R2_SB_n338), .C2(
        R2_SB_SB1_n629), .ZN(R2_SB_SB1_n632) );
  AOI221_X1 R2_SB_SB1_U202 ( .B1(R2_SB_SB1_n725), .B2(R2_SB_SB1_n728), .C1(
        R2_SB_SB1_n651), .C2(R2_SB_SB1_n789), .A(R2_SB_SB1_n632), .ZN(
        R2_SB_SB1_n643) );
  OAI222_X1 R2_SB_SB1_U201 ( .A1(R2_SB_SB1_n865), .A2(R2_SB_SB1_n785), .B1(
        R2_SB_SB1_n784), .B2(R2_SB_SB1_n905), .C1(R2_SB_SB1_n827), .C2(
        R2_SB_SB1_n897), .ZN(R2_SB_SB1_n786) );
  OAI211_X1 R2_SB_SB1_U200 ( .C1(R2_SB_SB1_n829), .C2(R2_SB_SB1_n770), .A(
        R2_SB_SB1_n769), .B(R2_SB_SB1_n768), .ZN(R2_SB_SB1_n788) );
  OAI211_X1 R2_SB_SB1_U199 ( .C1(R2_SB_SB1_n895), .C2(R2_SB_SB1_n848), .A(
        R2_SB_SB1_n777), .B(R2_SB_SB1_n887), .ZN(R2_SB_SB1_n787) );
  AOI221_X1 R2_SB_SB1_U198 ( .B1(R2_SB_SB1_n789), .B2(R2_SB_SB1_n788), .C1(
        R2_SB_n337), .C2(R2_SB_SB1_n787), .A(R2_SB_SB1_n786), .ZN(
        R2_SB_SB1_n823) );
  INV_X1 R2_SB_SB1_U197 ( .A(R2_SB_SB1_n656), .ZN(R2_SB_SB1_n859) );
  AOI211_X1 R2_SB_SB1_U196 ( .C1(R2_SB_SB1_n789), .C2(R2_SB_SB1_n812), .A(
        R2_SB_SB1_n882), .B(R2_SB_SB1_n727), .ZN(R2_SB_SB1_n577) );
  AOI211_X1 R2_SB_SB1_U195 ( .C1(R2_SB_SB1_n744), .C2(R2_SB_SB1_n843), .A(
        R2_SB_SB1_n730), .B(R2_SB_SB1_n792), .ZN(R2_SB_SB1_n509) );
  AOI21_X1 R2_SB_SB1_U194 ( .B1(R2_SB_SB1_n854), .B2(R2_SB_SB1_n881), .A(
        R2_SB_SB1_n767), .ZN(R2_SB_SB1_n477) );
  OAI222_X1 R2_SB_SB1_U193 ( .A1(R2_SB_SB1_n843), .A2(R2_SB_SB1_n885), .B1(
        R2_SB_SB1_n477), .B2(R2_SB_SB1_n845), .C1(R2_SB_SB1_n864), .C2(
        R2_SB_SB1_n878), .ZN(R2_SB_SB1_n479) );
  OAI22_X1 R2_SB_SB1_U192 ( .A1(R2_SB_SB1_n849), .A2(R2_SB_SB1_n648), .B1(
        R2_SB_SB1_n862), .B2(R2_SB_SB1_n844), .ZN(R2_SB_SB1_n478) );
  AOI211_X1 R2_SB_SB1_U191 ( .C1(R2_SB_SB1_n791), .C2(R2_SB_SB1_n812), .A(
        R2_SB_SB1_n479), .B(R2_SB_SB1_n478), .ZN(R2_SB_SB1_n480) );
  NOR3_X1 R2_SB_SB1_U190 ( .A1(R2_SB_SB1_n838), .A2(R2_SB_n337), .A3(
        R2_SB_SB1_n864), .ZN(R2_SB_SB1_n610) );
  AOI21_X1 R2_SB_SB1_U189 ( .B1(R2_SB_SB1_n858), .B2(R2_SB_SB1_n608), .A(
        R2_SB_SB1_n827), .ZN(R2_SB_SB1_n609) );
  AOI211_X1 R2_SB_SB1_U188 ( .C1(R2_SB_SB1_n646), .C2(R2_SB_SB1_n781), .A(
        R2_SB_SB1_n610), .B(R2_SB_SB1_n609), .ZN(R2_SB_SB1_n611) );
  INV_X1 R2_SB_SB1_U187 ( .A(R2_SB_SB1_n752), .ZN(R2_SB_SB1_n878) );
  NOR2_X1 R2_SB_SB1_U186 ( .A1(R2_SB_SB1_n857), .A2(R2_SB_SB1_n863), .ZN(
        R2_SB_SB1_n670) );
  INV_X1 R2_SB_SB1_U185 ( .A(R2_SB_SB1_n772), .ZN(R2_SB_SB1_n883) );
  INV_X1 R2_SB_SB1_U184 ( .A(R2_SB_SB1_n618), .ZN(R2_SB_SB1_n864) );
  OAI21_X1 R2_SB_SB1_U183 ( .B1(R2_SB_SB1_n856), .B2(R2_SB_SB1_n874), .A(
        R2_SB_SB1_n893), .ZN(R2_SB_SB1_n516) );
  AOI21_X1 R2_SB_SB1_U182 ( .B1(R2_SB_SB1_n781), .B2(R2_SB_SB1_n516), .A(
        R2_SB_SB1_n515), .ZN(R2_SB_SB1_n517) );
  AOI21_X1 R2_SB_SB1_U181 ( .B1(R2_SB_SB1_n900), .B2(R2_SB_SB1_n603), .A(
        R2_SB_SB1_n783), .ZN(R2_SB_SB1_n518) );
  OAI221_X1 R2_SB_SB1_U180 ( .B1(R2_SB_SB1_n518), .B2(R2_SB_SB1_n453), .C1(
        R2_SB_SB1_n838), .C2(R2_SB_SB1_n904), .A(R2_SB_SB1_n517), .ZN(
        R2_SB_SB1_n523) );
  AOI21_X1 R2_SB_SB1_U179 ( .B1(R2_SB_SB1_n646), .B2(R2_SB_SB1_n634), .A(
        R2_SB_SB1_n633), .ZN(R2_SB_SB1_n636) );
  OAI21_X1 R2_SB_SB1_U178 ( .B1(R2_SB_SB1_n747), .B2(R2_SB_SB1_n799), .A(
        R2_SB_SB1_n882), .ZN(R2_SB_SB1_n635) );
  NAND2_X1 R2_SB_SB1_U177 ( .A1(R2_SB_SB1_n828), .A2(R2_SB_SB1_n843), .ZN(
        R2_SB_SB1_n637) );
  OAI221_X1 R2_SB_SB1_U176 ( .B1(R2_SB_SB1_n910), .B2(R2_SB_SB1_n637), .C1(
        R2_SB_SB1_n636), .C2(R2_SB_SB1_n829), .A(R2_SB_SB1_n635), .ZN(
        R2_SB_SB1_n641) );
  OAI22_X1 R2_SB_SB1_U175 ( .A1(R2_SB_SB1_n857), .A2(R2_SB_SB1_n838), .B1(
        R2_SB_SB1_n832), .B2(R2_SB_SB1_n865), .ZN(R2_SB_SB1_n469) );
  OAI21_X1 R2_SB_SB1_U174 ( .B1(R2_SB_n338), .B2(R2_SB_SB1_n845), .A(
        R2_SB_SB1_n849), .ZN(R2_SB_SB1_n471) );
  AOI221_X1 R2_SB_SB1_U173 ( .B1(R2_SB_SB1_n744), .B2(R2_SB_SB1_n471), .C1(
        R2_SB_SB1_n470), .C2(R2_SB_SB1_n863), .A(R2_SB_SB1_n469), .ZN(
        R2_SB_SB1_n476) );
  AOI221_X1 R2_SB_SB1_U172 ( .B1(R2_SB_SB1_n882), .B2(R2_SB_SB1_n792), .C1(
        R2_SB_SB1_n627), .C2(R2_SB_SB1_n702), .A(R2_SB_SB1_n698), .ZN(
        R2_SB_SB1_n583) );
  NOR2_X1 R2_SB_SB1_U171 ( .A1(R2_SB_SB1_n813), .A2(R2_SB_SB1_n694), .ZN(
        R2_SB_SB1_n695) );
  OAI221_X1 R2_SB_SB1_U170 ( .B1(R2_SB_SB1_n695), .B2(R2_SB_SB1_n851), .C1(
        R2_SB_SB1_n856), .C2(R2_SB_SB1_n878), .A(R2_SB_SB1_n904), .ZN(
        R2_SB_SB1_n697) );
  INV_X1 R2_SB_SB1_U169 ( .A(R2_SB_SB1_n801), .ZN(R2_SB_SB1_n873) );
  AOI222_X1 R2_SB_SB1_U168 ( .A1(R2_SB_SB1_n771), .A2(R2_SB_SB1_n698), .B1(
        R2_SB_SB1_n781), .B2(R2_SB_SB1_n697), .C1(R2_SB_SB1_n696), .C2(
        R2_SB_SB1_n873), .ZN(R2_SB_SB1_n741) );
  AOI22_X1 R2_SB_SB1_U167 ( .A1(R2_SB_SB1_n758), .A2(R2_SB_SB1_n694), .B1(
        R2_SB_SB1_n779), .B2(R2_SB_SB1_n863), .ZN(R2_SB_SB1_n619) );
  OAI222_X1 R2_SB_SB1_U166 ( .A1(R2_SB_SB1_n864), .A2(R2_SB_SB1_n833), .B1(
        R2_SB_n337), .B2(R2_SB_SB1_n619), .C1(R2_SB_SB1_n858), .C2(
        R2_SB_SB1_n839), .ZN(R2_SB_SB1_n620) );
  AOI221_X1 R2_SB_SB1_U165 ( .B1(R2_SB_SB1_n789), .B2(R2_SB_SB1_n628), .C1(
        R2_SB_SB1_n778), .C2(R2_SB_SB1_n771), .A(R2_SB_SB1_n620), .ZN(
        R2_SB_SB1_n621) );
  NAND2_X1 R2_SB_SB1_U164 ( .A1(R2_SB_SB1_n848), .A2(R2_SB_SB1_n841), .ZN(
        R2_SB_SB1_n616) );
  INV_X1 R2_SB_SB1_U163 ( .A(R2_SB_SB1_n615), .ZN(R2_SB_SB1_n861) );
  AOI221_X1 R2_SB_SB1_U162 ( .B1(R2_SB_SB1_n747), .B2(R2_SB_SB1_n618), .C1(
        R2_SB_SB1_n617), .C2(R2_SB_SB1_n616), .A(R2_SB_SB1_n861), .ZN(
        R2_SB_SB1_n622) );
  OAI221_X1 R2_SB_SB1_U161 ( .B1(R2_SB_SB1_n870), .B2(R2_SB_SB1_n838), .C1(
        R2_SB_SB1_n840), .C2(R2_SB_SB1_n868), .A(R2_SB_SB1_n496), .ZN(
        R2_SB_SB1_n497) );
  OAI211_X1 R2_SB_SB1_U160 ( .C1(R2_SB_SB1_n879), .C2(R2_SB_SB1_n844), .A(
        R2_SB_SB1_n711), .B(R2_SB_SB1_n491), .ZN(R2_SB_SB1_n499) );
  AOI222_X1 R2_SB_SB1_U159 ( .A1(R2_SB_SB1_n499), .A2(R2_SB_SB1_n453), .B1(
        R2_SB_SB1_n498), .B2(R2_SB_SB1_n854), .C1(R2_SB_SB1_n752), .C2(
        R2_SB_SB1_n497), .ZN(R2_SB_SB1_n527) );
  OAI222_X1 R2_SB_SB1_U158 ( .A1(R2_SB_SB1_n865), .A2(R2_SB_SB1_n838), .B1(
        R2_SB_SB1_n699), .B2(R2_SB_SB1_n868), .C1(R2_SB_n338), .C2(
        R2_SB_SB1_n858), .ZN(R2_SB_SB1_n704) );
  OAI22_X1 R2_SB_SB1_U157 ( .A1(R2_SB_SB1_n864), .A2(R2_SB_SB1_n839), .B1(
        R2_SB_SB1_n700), .B2(R2_SB_SB1_n833), .ZN(R2_SB_SB1_n701) );
  AOI222_X1 R2_SB_SB1_U156 ( .A1(R2_SB_SB1_n772), .A2(R2_SB_SB1_n704), .B1(
        R2_SB_SB1_n882), .B2(R2_SB_SB1_n703), .C1(R2_SB_SB1_n702), .C2(
        R2_SB_SB1_n701), .ZN(R2_SB_SB1_n740) );
  NOR2_X1 R2_SB_SB1_U155 ( .A1(R2_SB_SB1_n881), .A2(R2_SB_SB1_n863), .ZN(
        R2_SB_SB1_n634) );
  OAI222_X1 R2_SB_SB1_U154 ( .A1(R2_SB_n338), .A2(R2_SB_SB1_n875), .B1(
        R2_SB_SB1_n883), .B2(R2_SB_SB1_n826), .C1(R2_SB_SB1_n905), .C2(
        R2_SB_SB1_n831), .ZN(R2_SB_SB1_n707) );
  AOI211_X1 R2_SB_SB1_U153 ( .C1(R2_SB_SB1_n709), .C2(R2_SB_SB1_n708), .A(
        R2_SB_SB1_n707), .B(R2_SB_SB1_n706), .ZN(R2_SB_SB1_n710) );
  OAI222_X1 R2_SB_SB1_U152 ( .A1(R2_SB_SB1_n833), .A2(R2_SB_SB1_n898), .B1(
        R2_SB_SB1_n710), .B2(R2_SB_SB1_n859), .C1(R2_SB_SB1_n832), .C2(
        R2_SB_SB1_n800), .ZN(R2_SB_SB1_n712) );
  INV_X1 R2_SB_SB1_U151 ( .A(R2_SB_SB1_n792), .ZN(R2_SB_SB1_n845) );
  OAI221_X1 R2_SB_SB1_U150 ( .B1(R2_SB_SB1_n833), .B2(R2_SB_SB1_n774), .C1(
        R2_SB_SB1_n509), .C2(R2_SB_SB1_n829), .A(R2_SB_SB1_n508), .ZN(
        R2_SB_SB1_n510) );
  AOI221_X1 R2_SB_SB1_U149 ( .B1(R2_SB_SB1_n507), .B2(R2_SB_SB1_n506), .C1(
        R2_SB_SB1_n780), .C2(R2_SB_SB1_n684), .A(R2_SB_SB1_n505), .ZN(
        R2_SB_SB1_n512) );
  AOI221_X1 R2_SB_SB1_U148 ( .B1(R2_SB_SB1_n743), .B2(R2_SB_SB1_n684), .C1(
        R2_SB_SB1_n780), .C2(R2_SB_SB1_n627), .A(R2_SB_SB1_n510), .ZN(
        R2_SB_SB1_n511) );
  OAI222_X1 R2_SB_SB1_U147 ( .A1(R2_SB_SB1_n512), .A2(R2_SB_SB1_n905), .B1(
        R2_SB_SB1_n511), .B2(R2_SB_SB1_n883), .C1(R2_SB_SB1_n884), .C2(
        R2_SB_SB1_n844), .ZN(R2_SB_SB1_n513) );
  INV_X1 R2_SB_SB1_U146 ( .A(R2_SB_SB1_n659), .ZN(R2_SB_SB1_n867) );
  AOI221_X1 R2_SB_SB1_U145 ( .B1(R2_SB_SB1_n794), .B2(R2_SB_SB1_n730), .C1(
        R2_SB_SB1_n742), .C2(R2_SB_SB1_n780), .A(R2_SB_SB1_n867), .ZN(
        R2_SB_SB1_n574) );
  NOR4_X1 R2_SB_SB1_U144 ( .A1(R2_SB_SB1_n452), .A2(R2_SB_SB1_n872), .A3(
        R2_SB_SB1_n849), .A4(R2_SB_SB1_n862), .ZN(R2_SB_SB1_n640) );
  NOR2_X1 R2_SB_SB1_U143 ( .A1(R2_SB_SB1_n89), .A2(R2_SB_SB1_n843), .ZN(
        R2_SB_SB1_n603) );
  NOR2_X1 R2_SB_SB1_U142 ( .A1(R2_SB_SB1_n872), .A2(R2_SB_SB1_n863), .ZN(
        R2_SB_SB1_n812) );
  NOR2_X1 R2_SB_SB1_U141 ( .A1(R2_SB_SB1_n863), .A2(R2_SB_SB1_n854), .ZN(
        R2_SB_SB1_n507) );
  AOI222_X1 R2_SB_SB1_U140 ( .A1(R2_SB_SB1_n782), .A2(R2_SB_SB1_n781), .B1(
        R2_SB_SB1_n780), .B2(R2_SB_SB1_n779), .C1(R2_SB_SB1_n778), .C2(
        R2_SB_SB1_n791), .ZN(R2_SB_SB1_n784) );
  INV_X1 R2_SB_SB1_U139 ( .A(R2_SB_SB1_n795), .ZN(R2_SB_SB1_n838) );
  AOI22_X1 R2_SB_SB1_U138 ( .A1(R2_SB_SB1_n724), .A2(R2_SB_SB1_n810), .B1(
        R2_SB_SB1_n744), .B2(R2_SB_SB1_n723), .ZN(R2_SB_SB1_n726) );
  INV_X1 R2_SB_SB1_U137 ( .A(R2_SB_SB1_n722), .ZN(R2_SB_SB1_n896) );
  INV_X1 R2_SB_SB1_U136 ( .A(R2_SB_SB1_n725), .ZN(R2_SB_SB1_n846) );
  OAI222_X1 R2_SB_SB1_U135 ( .A1(R2_SB_SB1_n849), .A2(R2_SB_SB1_n896), .B1(
        R2_SB_SB1_n726), .B2(R2_SB_SB1_n878), .C1(R2_SB_SB1_n846), .C2(
        R2_SB_SB1_n910), .ZN(R2_SB_SB1_n735) );
  OAI222_X1 R2_SB_SB1_U134 ( .A1(R2_SB_SB1_n853), .A2(R2_SB_SB1_n829), .B1(
        R2_SB_SB1_n608), .B2(R2_SB_SB1_n826), .C1(R2_SB_SB1_n870), .C2(
        R2_SB_SB1_n831), .ZN(R2_SB_SB1_n465) );
  NOR3_X1 R2_SB_SB1_U133 ( .A1(R2_SB_SB1_n877), .A2(R2_SB_SB1_n638), .A3(
        R2_SB_SB1_n679), .ZN(R2_SB_SB1_n466) );
  INV_X1 R2_SB_SB1_U132 ( .A(R2_SB_SB1_n465), .ZN(R2_SB_SB1_n871) );
  OAI222_X1 R2_SB_SB1_U131 ( .A1(R2_SB_SB1_n871), .A2(R2_SB_SB1_n883), .B1(
        R2_SB_SB1_n849), .B2(R2_SB_SB1_n769), .C1(R2_SB_SB1_n466), .C2(
        R2_SB_SB1_n834), .ZN(R2_SB_SB1_n484) );
  INV_X1 R2_SB_SB1_U130 ( .A(R2_SB_SB1_n782), .ZN(R2_SB_SB1_n849) );
  NOR2_X1 R2_SB_SB1_U129 ( .A1(R2_SB_SB1_n830), .A2(R2_SB_SB1_n854), .ZN(
        R2_SB_SB1_n627) );
  NOR2_X1 R2_SB_SB1_U128 ( .A1(R2_SB_SB1_n881), .A2(R2_SB_SB1_n872), .ZN(
        R2_SB_SB1_n669) );
  INV_X1 R2_SB_SB1_U127 ( .A(R2_SB_SB1_n702), .ZN(R2_SB_SB1_n905) );
  NOR2_X1 R2_SB_SB1_U126 ( .A1(R2_SB_SB1_n453), .A2(R2_SB_SB1_n830), .ZN(
        R2_SB_SB1_n766) );
  NOR3_X1 R2_SB_SB1_U125 ( .A1(R2_SB_SB1_n828), .A2(R2_SB_SB1_n854), .A3(
        R2_SB_SB1_n908), .ZN(R2_SB_SB1_n673) );
  NOR2_X1 R2_SB_SB1_U124 ( .A1(R2_SB_SB1_n89), .A2(R2_SB_SB1_n830), .ZN(
        R2_SB_SB1_n771) );
  NOR2_X1 R2_SB_SB1_U123 ( .A1(R2_SB_SB1_n863), .A2(R2_SB_SB1_n843), .ZN(
        R2_SB_SB1_n778) );
  NOR2_X1 R2_SB_SB1_U122 ( .A1(R2_SB_SB1_n830), .A2(R2_SB_n338), .ZN(
        R2_SB_SB1_n779) );
  AOI21_X1 R2_SB_SB1_U121 ( .B1(R2_SB_SB1_n826), .B2(R2_SB_SB1_n833), .A(
        R2_SB_SB1_n800), .ZN(R2_SB_SB1_n549) );
  INV_X1 R2_SB_SB1_U120 ( .A(R2_SB_SB1_n549), .ZN(R2_SB_SB1_n902) );
  AND3_X1 R2_SB_SB1_U119 ( .A1(R2_SB_SB1_n548), .A2(R2_SB_SB1_n838), .A3(
        R2_SB_SB1_n849), .ZN(R2_SB_SB1_n550) );
  OR3_X1 R2_SB_SB1_U118 ( .A1(R2_SB_SB1_n864), .A2(R2_SB_SB1_n814), .A3(
        R2_SB_SB1_n890), .ZN(R2_SB_SB1_n815) );
  INV_X1 R2_SB_SB1_U117 ( .A(R2_SB_SB1_n519), .ZN(R2_SB_SB1_n886) );
  INV_X1 R2_SB_SB1_U116 ( .A(R2_SB_SB1_n790), .ZN(R2_SB_SB1_n866) );
  NAND2_X1 R2_SB_SB1_U115 ( .A1(R2_SB_SB1_n874), .A2(R2_SB_SB1_n901), .ZN(
        R2_SB_SB1_n728) );
  NAND2_X1 R2_SB_SB1_U114 ( .A1(R2_SB_SB1_n890), .A2(R2_SB_SB1_n874), .ZN(
        R2_SB_SB1_n536) );
  NAND2_X1 R2_SB_SB1_U113 ( .A1(R2_SB_SB1_n836), .A2(R2_SB_SB1_n826), .ZN(
        R2_SB_SB1_n723) );
  NAND2_X1 R2_SB_SB1_U112 ( .A1(R2_SB_SB1_n905), .A2(R2_SB_SB1_n875), .ZN(
        R2_SB_SB1_n589) );
  INV_X1 R2_SB_SB1_U111 ( .A(R2_SB_SB1_n627), .ZN(R2_SB_SB1_n856) );
  NAND2_X1 R2_SB_SB1_U110 ( .A1(R2_SB_SB1_n836), .A2(R2_SB_SB1_n829), .ZN(
        R2_SB_SB1_n748) );
  AND2_X1 R2_SB_SB1_U109 ( .A1(R2_SB_SB1_n766), .A2(R2_SB_SB1_n671), .ZN(
        R2_SB_SB1_n555) );
  INV_X1 R2_SB_SB1_U108 ( .A(R2_SB_SB1_n812), .ZN(R2_SB_SB1_n875) );
  OAI21_X1 R2_SB_SB1_U107 ( .B1(R2_SB_SB1_n847), .B2(R2_SB_SB1_n895), .A(
        R2_SB_SB1_n800), .ZN(R2_SB_SB1_n806) );
  NAND2_X1 R2_SB_SB1_U106 ( .A1(R2_SB_SB1_n628), .A2(R2_SB_SB1_n634), .ZN(
        R2_SB_SB1_n769) );
  NAND2_X1 R2_SB_SB1_U105 ( .A1(R2_SB_SB1_n507), .A2(R2_SB_SB1_n669), .ZN(
        R2_SB_SB1_n588) );
  INV_X1 R2_SB_SB1_U104 ( .A(R2_SB_SB1_n634), .ZN(R2_SB_SB1_n903) );
  INV_X1 R2_SB_SB1_U103 ( .A(R2_SB_SB1_n778), .ZN(R2_SB_SB1_n865) );
  NOR2_X1 R2_SB_SB1_U102 ( .A1(R2_SB_SB1_n730), .A2(R2_SB_SB1_n758), .ZN(
        R2_SB_SB1_n685) );
  AOI21_X1 R2_SB_SB1_U101 ( .B1(R2_SB_SB1_n588), .B2(R2_SB_SB1_n773), .A(
        R2_SB_SB1_n836), .ZN(R2_SB_SB1_n460) );
  AOI21_X1 R2_SB_SB1_U100 ( .B1(R2_SB_SB1_n802), .B2(R2_SB_SB1_n801), .A(
        R2_SB_SB1_n835), .ZN(R2_SB_SB1_n803) );
  INV_X1 R2_SB_SB1_U99 ( .A(R2_SB_SB1_n672), .ZN(R2_SB_SB1_n888) );
  NOR4_X1 R2_SB_SB1_U98 ( .A1(R2_SB_SB1_n675), .A2(R2_SB_SB1_n888), .A3(
        R2_SB_SB1_n674), .A4(R2_SB_SB1_n673), .ZN(R2_SB_SB1_n676) );
  NAND2_X1 R2_SB_SB1_U97 ( .A1(R2_SB_SB1_n778), .A2(R2_SB_SB1_n669), .ZN(
        R2_SB_SB1_n573) );
  INV_X1 R2_SB_SB1_U96 ( .A(R2_SB_SB1_n648), .ZN(R2_SB_SB1_n882) );
  NOR2_X1 R2_SB_SB1_U95 ( .A1(R2_SB_SB1_n849), .A2(R2_SB_SB1_n89), .ZN(
        R2_SB_SB1_n502) );
  NOR2_X1 R2_SB_SB1_U94 ( .A1(R2_SB_SB1_n851), .A2(R2_SB_n338), .ZN(
        R2_SB_SB1_n470) );
  NOR2_X1 R2_SB_SB1_U93 ( .A1(R2_SB_SB1_n853), .A2(R2_SB_SB1_n903), .ZN(
        R2_SB_SB1_n514) );
  INV_X1 R2_SB_SB1_U92 ( .A(R2_SB_SB1_n604), .ZN(R2_SB_SB1_n844) );
  NOR2_X1 R2_SB_SB1_U91 ( .A1(R2_SB_SB1_n862), .A2(R2_SB_SB1_n883), .ZN(
        R2_SB_SB1_n534) );
  INV_X1 R2_SB_SB1_U90 ( .A(R2_SB_SB1_n603), .ZN(R2_SB_SB1_n848) );
  INV_X1 R2_SB_SB1_U89 ( .A(R2_SB_SB1_n802), .ZN(R2_SB_SB1_n877) );
  NOR2_X1 R2_SB_SB1_U88 ( .A1(R2_SB_SB1_n905), .A2(R2_SB_SB1_n866), .ZN(
        R2_SB_SB1_n671) );
  OAI22_X1 R2_SB_SB1_U87 ( .A1(R2_SB_SB1_n730), .A2(R2_SB_SB1_n905), .B1(
        R2_SB_SB1_n901), .B2(R2_SB_SB1_n851), .ZN(R2_SB_SB1_n462) );
  OAI22_X1 R2_SB_SB1_U86 ( .A1(R2_SB_SB1_n875), .A2(R2_SB_SB1_n833), .B1(
        R2_SB_SB1_n874), .B2(R2_SB_SB1_n832), .ZN(R2_SB_SB1_n804) );
  OAI22_X1 R2_SB_SB1_U85 ( .A1(R2_SB_SB1_n665), .A2(R2_SB_SB1_n892), .B1(
        R2_SB_SB1_n841), .B2(R2_SB_SB1_n801), .ZN(R2_SB_SB1_n666) );
  INV_X1 R2_SB_SB1_U84 ( .A(R2_SB_SB1_n758), .ZN(R2_SB_SB1_n847) );
  AOI21_X1 R2_SB_SB1_U83 ( .B1(R2_SB_SB1_n868), .B2(R2_SB_SB1_n845), .A(
        R2_SB_SB1_n785), .ZN(R2_SB_SB1_n687) );
  OAI22_X1 R2_SB_SB1_U82 ( .A1(R2_SB_SB1_n831), .A2(R2_SB_SB1_n895), .B1(
        R2_SB_n337), .B2(R2_SB_SB1_n648), .ZN(R2_SB_SB1_n532) );
  AOI22_X1 R2_SB_SB1_U81 ( .A1(R2_SB_SB1_n758), .A2(R2_SB_n338), .B1(
        R2_SB_SB1_n771), .B2(R2_SB_SB1_n452), .ZN(R2_SB_SB1_n699) );
  INV_X1 R2_SB_SB1_U80 ( .A(R2_SB_SB1_n771), .ZN(R2_SB_SB1_n831) );
  NOR2_X1 R2_SB_SB1_U79 ( .A1(R2_SB_SB1_n842), .A2(R2_SB_SB1_n898), .ZN(
        R2_SB_SB1_n675) );
  NOR2_X1 R2_SB_SB1_U78 ( .A1(R2_SB_SB1_n868), .A2(R2_SB_SB1_n890), .ZN(
        R2_SB_SB1_n576) );
  NOR2_X1 R2_SB_SB1_U77 ( .A1(R2_SB_SB1_n774), .A2(R2_SB_SB1_n890), .ZN(
        R2_SB_SB1_n565) );
  NOR2_X1 R2_SB_SB1_U76 ( .A1(R2_SB_SB1_n845), .A2(R2_SB_SB1_n89), .ZN(
        R2_SB_SB1_n725) );
  NOR2_X1 R2_SB_SB1_U75 ( .A1(R2_SB_SB1_n853), .A2(R2_SB_SB1_n890), .ZN(
        R2_SB_SB1_n633) );
  NOR2_X1 R2_SB_SB1_U74 ( .A1(R2_SB_SB1_n868), .A2(R2_SB_SB1_n905), .ZN(
        R2_SB_SB1_n754) );
  NOR2_X1 R2_SB_SB1_U73 ( .A1(R2_SB_SB1_n869), .A2(R2_SB_SB1_n905), .ZN(
        R2_SB_SB1_n698) );
  NOR2_X1 R2_SB_SB1_U72 ( .A1(R2_SB_SB1_n898), .A2(R2_SB_SB1_n845), .ZN(
        R2_SB_SB1_n756) );
  NOR2_X1 R2_SB_SB1_U71 ( .A1(R2_SB_SB1_n774), .A2(R2_SB_SB1_n905), .ZN(
        R2_SB_SB1_n638) );
  NOR2_X1 R2_SB_SB1_U70 ( .A1(R2_SB_SB1_n870), .A2(R2_SB_SB1_n890), .ZN(
        R2_SB_SB1_n727) );
  OAI22_X1 R2_SB_SB1_U69 ( .A1(R2_SB_SB1_n453), .A2(R2_SB_SB1_n879), .B1(
        R2_SB_SB1_n89), .B2(R2_SB_SB1_n880), .ZN(R2_SB_SB1_n538) );
  AOI211_X1 R2_SB_SB1_U68 ( .C1(R2_SB_SB1_n576), .C2(R2_SB_SB1_n89), .A(
        R2_SB_SB1_n538), .B(R2_SB_SB1_n722), .ZN(R2_SB_SB1_n543) );
  INV_X1 R2_SB_SB1_U67 ( .A(R2_SB_SB1_n779), .ZN(R2_SB_SB1_n833) );
  NOR3_X1 R2_SB_SB1_U66 ( .A1(R2_SB_SB1_n841), .A2(R2_SB_SB1_n858), .A3(
        R2_SB_SB1_n874), .ZN(R2_SB_SB1_n521) );
  INV_X1 R2_SB_SB1_U65 ( .A(R2_SB_SB1_n766), .ZN(R2_SB_SB1_n835) );
  NOR2_X1 R2_SB_SB1_U64 ( .A1(R2_SB_SB1_n838), .A2(R2_SB_SB1_n453), .ZN(
        R2_SB_SB1_n742) );
  INV_X1 R2_SB_SB1_U63 ( .A(R2_SB_SB1_n730), .ZN(R2_SB_SB1_n858) );
  NOR2_X1 R2_SB_SB1_U62 ( .A1(R2_SB_SB1_n878), .A2(R2_SB_SB1_n869), .ZN(
        R2_SB_SB1_n713) );
  NOR2_X1 R2_SB_SB1_U61 ( .A1(R2_SB_SB1_n833), .A2(R2_SB_SB1_n453), .ZN(
        R2_SB_SB1_n799) );
  AOI22_X1 R2_SB_SB1_U60 ( .A1(R2_SB_SB1_n877), .A2(R2_SB_SB1_n452), .B1(
        R2_SB_SB1_n781), .B2(R2_SB_SB1_n669), .ZN(R2_SB_SB1_n500) );
  OAI211_X1 R2_SB_SB1_U59 ( .C1(R2_SB_SB1_n89), .C2(R2_SB_SB1_n893), .A(
        R2_SB_SB1_n907), .B(R2_SB_SB1_n500), .ZN(R2_SB_SB1_n501) );
  AOI222_X1 R2_SB_SB1_U58 ( .A1(R2_SB_SB1_n591), .A2(R2_SB_SB1_n748), .B1(
        R2_SB_SB1_n502), .B2(R2_SB_SB1_n679), .C1(R2_SB_SB1_n758), .C2(
        R2_SB_SB1_n501), .ZN(R2_SB_SB1_n526) );
  OAI222_X1 R2_SB_SB1_U57 ( .A1(R2_SB_SB1_n845), .A2(R2_SB_SB1_n880), .B1(
        R2_SB_SB1_n835), .B2(R2_SB_SB1_n898), .C1(R2_SB_SB1_n836), .C2(
        R2_SB_SB1_n894), .ZN(R2_SB_SB1_n602) );
  NOR2_X1 R2_SB_SB1_U56 ( .A1(R2_SB_SB1_n883), .A2(R2_SB_SB1_n869), .ZN(
        R2_SB_SB1_n755) );
  NOR2_X1 R2_SB_SB1_U55 ( .A1(R2_SB_SB1_n862), .A2(R2_SB_SB1_n890), .ZN(
        R2_SB_SB1_n753) );
  NOR2_X1 R2_SB_SB1_U54 ( .A1(R2_SB_SB1_n862), .A2(R2_SB_SB1_n905), .ZN(
        R2_SB_SB1_n759) );
  NOR2_X1 R2_SB_SB1_U53 ( .A1(R2_SB_SB1_n862), .A2(R2_SB_SB1_n878), .ZN(
        R2_SB_SB1_n591) );
  NOR2_X1 R2_SB_SB1_U52 ( .A1(R2_SB_SB1_n869), .A2(R2_SB_SB1_n890), .ZN(
        R2_SB_SB1_n679) );
  INV_X1 R2_SB_SB1_U51 ( .A(R2_SB_SB1_n669), .ZN(R2_SB_SB1_n890) );
  NOR2_X2 R2_SB_SB1_U50 ( .A1(R2_SB_SB1_n89), .A2(R2_SB_SB1_n453), .ZN(
        R2_SB_SB1_n781) );
  NOR2_X2 R2_SB_SB1_U49 ( .A1(R2_SB_SB1_n89), .A2(R2_SB_SB1_n452), .ZN(
        R2_SB_SB1_n684) );
  NOR3_X1 R2_SB_SB1_U48 ( .A1(R2_SB_SB1_n878), .A2(R2_SB_SB1_n866), .A3(
        R2_SB_SB1_n838), .ZN(R2_SB_SB1_n674) );
  NOR2_X1 R2_SB_SB1_U47 ( .A1(R2_SB_SB1_n840), .A2(R2_SB_SB1_n452), .ZN(
        R2_SB_SB1_n747) );
  NOR2_X1 R2_SB_SB1_U46 ( .A1(R2_SB_SB1_n453), .A2(R2_SB_n338), .ZN(
        R2_SB_SB1_n810) );
  INV_X1 R2_SB_SB1_U45 ( .A(R2_SB_SB1_n633), .ZN(R2_SB_SB1_n891) );
  INV_X1 R2_SB_SB1_U44 ( .A(R2_SB_SB1_n534), .ZN(R2_SB_SB1_n885) );
  INV_X1 R2_SB_SB1_U43 ( .A(R2_SB_SB1_n470), .ZN(R2_SB_SB1_n852) );
  INV_X1 R2_SB_SB1_U42 ( .A(R2_SB_SB1_n502), .ZN(R2_SB_SB1_n850) );
  INV_X1 R2_SB_SB1_U41 ( .A(R2_SB_SB1_n514), .ZN(R2_SB_SB1_n904) );
  INV_X1 R2_SB_SB1_U40 ( .A(R2_SB_SB1_n698), .ZN(R2_SB_SB1_n906) );
  INV_X1 R2_SB_SB1_U39 ( .A(R2_SB_SB1_n638), .ZN(R2_SB_SB1_n908) );
  INV_X1 R2_SB_SB1_U38 ( .A(R2_SB_SB1_n565), .ZN(R2_SB_SB1_n892) );
  INV_X1 R2_SB_SB1_U37 ( .A(R2_SB_SB1_n753), .ZN(R2_SB_SB1_n893) );
  INV_X1 R2_SB_SB1_U36 ( .A(R2_SB_SB1_n727), .ZN(R2_SB_SB1_n894) );
  INV_X1 R2_SB_SB1_U35 ( .A(R2_SB_SB1_n755), .ZN(R2_SB_SB1_n884) );
  INV_X1 R2_SB_SB1_U34 ( .A(R2_SB_SB1_n799), .ZN(R2_SB_SB1_n834) );
  NAND2_X1 R2_SB_SB1_U33 ( .A1(R2_SB_SB1_n781), .A2(R2_SB_SB1_n671), .ZN(
        R2_SB_SB1_n716) );
  INV_X1 R2_SB_SB1_U32 ( .A(R2_SB_SB1_n588), .ZN(R2_SB_SB1_n900) );
  INV_X1 R2_SB_SB1_U31 ( .A(R2_SB_SB1_n759), .ZN(R2_SB_SB1_n907) );
  INV_X1 R2_SB_SB1_U30 ( .A(R2_SB_SB1_n747), .ZN(R2_SB_SB1_n841) );
  INV_X1 R2_SB_SB1_U29 ( .A(R2_SB_SB1_n713), .ZN(R2_SB_SB1_n879) );
  INV_X1 R2_SB_SB1_U28 ( .A(R2_SB_SB1_n591), .ZN(R2_SB_SB1_n880) );
  INV_X1 R2_SB_SB1_U27 ( .A(R2_SB_SB1_n742), .ZN(R2_SB_SB1_n839) );
  AOI21_X1 R2_SB_SB1_U26 ( .B1(R2_SB_SB1_n848), .B2(R2_SB_SB1_n852), .A(
        R2_SB_SB1_n910), .ZN(R2_SB_SB1_n461) );
  AOI21_X1 R2_SB_SB1_U25 ( .B1(R2_SB_SB1_n831), .B2(R2_SB_SB1_n835), .A(
        R2_SB_SB1_n890), .ZN(R2_SB_SB1_n796) );
  INV_X1 R2_SB_SB1_U24 ( .A(R2_SB_SB1_n684), .ZN(R2_SB_SB1_n827) );
  AOI22_X1 R2_SB_SB1_U23 ( .A1(R2_SB_SB1_n877), .A2(R2_SB_n338), .B1(
        R2_SB_SB1_n713), .B2(R2_SB_SB1_n828), .ZN(R2_SB_SB1_n649) );
  INV_X1 R2_SB_SB1_U22 ( .A(R2_SB_SB1_n754), .ZN(R2_SB_SB1_n910) );
  INV_X1 R2_SB_SB1_U21 ( .A(R2_SB_SB1_n781), .ZN(R2_SB_SB1_n828) );
  INV_X1 R2_SB_SB1_U20 ( .A(R2_SB_SB1_n576), .ZN(R2_SB_SB1_n898) );
  INV_X1 R2_SB_SB1_U19 ( .A(R2_SB_SB1_n679), .ZN(R2_SB_SB1_n895) );
  NOR2_X1 R2_SB_SB1_U18 ( .A1(R2_SB_SB1_n831), .A2(R2_SB_SB1_n452), .ZN(
        R2_SB_SB1_n708) );
  OAI221_X1 R2_SB_SB1_U17 ( .B1(R2_SB_n338), .B2(R2_SB_SB1_n906), .C1(
        R2_SB_SB1_n890), .C2(R2_SB_SB1_n826), .A(R2_SB_SB1_n769), .ZN(
        R2_SB_SB1_n590) );
  NOR2_X1 R2_SB_SB1_U16 ( .A1(R2_SB_SB1_n895), .A2(R2_SB_SB1_n452), .ZN(
        R2_SB_SB1_n722) );
  INV_X1 R2_SB_SB1_U15 ( .A(R2_SB_SB1_n810), .ZN(R2_SB_SB1_n829) );
  NOR2_X1 R2_SB_SB1_U14 ( .A1(R2_SB_n337), .A2(R2_SB_n338), .ZN(R2_SB_SB1_n628) );
  INV_X1 R2_SB_SB1_U13 ( .A(R2_SB_SB1_n708), .ZN(R2_SB_SB1_n832) );
  INV_X1 R2_SB_SB1_U12 ( .A(R2_SB_SB1_n628), .ZN(R2_SB_SB1_n826) );
  NOR2_X1 R2_SB_SB1_U11 ( .A1(R2_SB_SB1_n863), .A2(R2_SB_n341), .ZN(
        R2_SB_SB1_n744) );
  NOR2_X1 R2_SB_SB1_U10 ( .A1(R2_SB_SB1_n881), .A2(R2_SB_n343), .ZN(
        R2_SB_SB1_n772) );
  NOR2_X1 R2_SB_SB1_U9 ( .A1(R2_SB_SB1_n89), .A2(R2_SB_n339), .ZN(
        R2_SB_SB1_n791) );
  NOR2_X1 R2_SB_SB1_U8 ( .A1(R2_SB_SB1_n872), .A2(R2_SB_n344), .ZN(
        R2_SB_SB1_n752) );
  NOR2_X1 R2_SB_SB1_U7 ( .A1(R2_SB_SB1_n854), .A2(R2_SB_SB1_n843), .ZN(
        R2_SB_SB1_n730) );
  NOR2_X1 R2_SB_SB1_U6 ( .A1(R2_SB_SB1_n843), .A2(R2_SB_n342), .ZN(
        R2_SB_SB1_n780) );
  NOR2_X1 R2_SB_SB1_U5 ( .A1(R2_SB_n339), .A2(R2_SB_n340), .ZN(R2_SB_SB1_n743)
         );
  INV_X1 R2_SB_SB1_U4 ( .A(R2_SB_n340), .ZN(R2_SB_SB1_n843) );
  NOR2_X1 R2_SB_SB1_U3 ( .A1(R2_SB_SB1_n453), .A2(R2_SB_n339), .ZN(
        R2_SB_SB1_n696) );
  NOR2_X1 R2_SB_SB1_U2 ( .A1(R2_SB_SB1_n881), .A2(R2_SB_n342), .ZN(
        R2_SB_SB1_n798) );
  NOR2_X1 R2_SB_SB1_U1 ( .A1(R2_SB_SB1_n843), .A2(R2_SB_n341), .ZN(
        R2_SB_SB1_n789) );
  NAND3_X1 R2_SB_SB1_U464 ( .A1(R2_SB_SB1_n772), .A2(R2_SB_SB1_n670), .A3(
        R2_SB_SB1_n794), .ZN(R2_SB_SB1_n519) );
  OAI33_X1 R2_SB_SB1_U463 ( .A1(R2_SB_SB1_n838), .A2(R2_SB_SB1_n858), .A3(
        R2_SB_SB1_n905), .B1(R2_SB_SB1_n853), .B2(R2_SB_SB1_n830), .B3(
        R2_SB_SB1_n874), .ZN(R2_SB_SB1_n467) );
  NAND3_X1 R2_SB_SB1_U462 ( .A1(R2_SB_SB1_n507), .A2(R2_SB_SB1_n702), .A3(
        R2_SB_SB1_n758), .ZN(R2_SB_SB1_n677) );
  OAI33_X1 R2_SB_SB1_U461 ( .A1(R2_SB_SB1_n828), .A2(R2_SB_n344), .A3(
        R2_SB_n339), .B1(R2_SB_SB1_n472), .B2(R2_SB_SB1_n854), .B3(
        R2_SB_SB1_n829), .ZN(R2_SB_SB1_n473) );
  NAND4_X1 R2_SB_SB1_U460 ( .A1(R2_SB_SB1_n488), .A2(R2_SB_SB1_n487), .A3(
        R2_SB_SB1_n486), .A4(R2_SB_SB1_n485), .ZN(R2_SB_n329) );
  NAND3_X1 R2_SB_SB1_U459 ( .A1(R2_SB_SB1_n781), .A2(R2_SB_n339), .A3(
        R2_SB_SB1_n798), .ZN(R2_SB_SB1_n494) );
  NAND4_X1 R2_SB_SB1_U458 ( .A1(R2_SB_SB1_n743), .A2(R2_SB_SB1_n628), .A3(
        R2_SB_SB1_n767), .A4(R2_SB_n344), .ZN(R2_SB_SB1_n493) );
  NAND3_X1 R2_SB_SB1_U457 ( .A1(R2_SB_SB1_n813), .A2(R2_SB_SB1_n830), .A3(
        R2_SB_SB1_n684), .ZN(R2_SB_SB1_n492) );
  NAND3_X1 R2_SB_SB1_U456 ( .A1(R2_SB_SB1_n494), .A2(R2_SB_SB1_n493), .A3(
        R2_SB_SB1_n492), .ZN(R2_SB_SB1_n498) );
  NAND3_X1 R2_SB_SB1_U455 ( .A1(R2_SB_SB1_n844), .A2(R2_SB_SB1_n836), .A3(
        R2_SB_SB1_n548), .ZN(R2_SB_SB1_n506) );
  OAI33_X1 R2_SB_SB1_U454 ( .A1(R2_SB_SB1_n827), .A2(R2_SB_SB1_n856), .A3(
        R2_SB_SB1_n903), .B1(R2_SB_SB1_n898), .B2(R2_SB_SB1_n843), .B3(
        R2_SB_SB1_n826), .ZN(R2_SB_SB1_n515) );
  NAND3_X1 R2_SB_SB1_U453 ( .A1(R2_SB_SB1_n671), .A2(R2_SB_SB1_n453), .A3(
        R2_SB_n339), .ZN(R2_SB_SB1_n816) );
  NAND3_X1 R2_SB_SB1_U452 ( .A1(R2_SB_SB1_n670), .A2(R2_SB_SB1_n669), .A3(
        R2_SB_SB1_n779), .ZN(R2_SB_SB1_n672) );
  NAND3_X1 R2_SB_SB1_U451 ( .A1(R2_SB_SB1_n816), .A2(R2_SB_SB1_n519), .A3(
        R2_SB_SB1_n672), .ZN(R2_SB_SB1_n522) );
  OAI33_X1 R2_SB_SB1_U450 ( .A1(R2_SB_SB1_n832), .A2(R2_SB_SB1_n864), .A3(
        R2_SB_SB1_n890), .B1(R2_SB_SB1_n829), .B2(R2_SB_n344), .B3(
        R2_SB_SB1_n866), .ZN(R2_SB_SB1_n520) );
  NAND4_X1 R2_SB_SB1_U449 ( .A1(R2_SB_SB1_n527), .A2(R2_SB_SB1_n526), .A3(
        R2_SB_SB1_n525), .A4(R2_SB_SB1_n524), .ZN(R2_SB_n330) );
  NAND3_X1 R2_SB_SB1_U448 ( .A1(R2_SB_SB1_n744), .A2(R2_SB_SB1_n603), .A3(
        R2_SB_SB1_n696), .ZN(R2_SB_SB1_n546) );
  NAND3_X1 R2_SB_SB1_U447 ( .A1(R2_SB_SB1_n684), .A2(R2_SB_SB1_n854), .A3(
        R2_SB_SB1_n709), .ZN(R2_SB_SB1_n582) );
  OAI33_X1 R2_SB_SB1_U446 ( .A1(R2_SB_SB1_n859), .A2(R2_SB_SB1_n830), .A3(
        R2_SB_SB1_n901), .B1(R2_SB_SB1_n876), .B2(R2_SB_n338), .B3(
        R2_SB_SB1_n685), .ZN(R2_SB_SB1_n557) );
  NAND4_X1 R2_SB_SB1_U445 ( .A1(R2_SB_SB1_n561), .A2(R2_SB_SB1_n560), .A3(
        R2_SB_SB1_n559), .A4(R2_SB_SB1_n558), .ZN(R2_SB_n331) );
  NAND3_X1 R2_SB_SB1_U444 ( .A1(R2_SB_SB1_n830), .A2(R2_SB_SB1_n872), .A3(
        R2_SB_SB1_n709), .ZN(R2_SB_SB1_n566) );
  NAND4_X1 R2_SB_SB1_U443 ( .A1(R2_SB_SB1_n566), .A2(R2_SB_SB1_n894), .A3(
        R2_SB_SB1_n800), .A4(R2_SB_SB1_n648), .ZN(R2_SB_SB1_n569) );
  NAND3_X1 R2_SB_SB1_U442 ( .A1(R2_SB_n337), .A2(R2_SB_n340), .A3(
        R2_SB_SB1_n744), .ZN(R2_SB_SB1_n659) );
  NAND3_X1 R2_SB_SB1_U441 ( .A1(R2_SB_SB1_n758), .A2(R2_SB_SB1_n854), .A3(
        R2_SB_SB1_n709), .ZN(R2_SB_SB1_n587) );
  NAND3_X1 R2_SB_SB1_U440 ( .A1(R2_SB_SB1_n743), .A2(R2_SB_n337), .A3(
        R2_SB_SB1_n882), .ZN(R2_SB_SB1_n592) );
  NAND4_X1 R2_SB_SB1_U439 ( .A1(R2_SB_SB1_n601), .A2(R2_SB_SB1_n600), .A3(
        R2_SB_SB1_n599), .A4(R2_SB_SB1_n598), .ZN(R2_SB_n332) );
  NAND4_X1 R2_SB_SB1_U438 ( .A1(R2_SB_SB1_n645), .A2(R2_SB_SB1_n644), .A3(
        R2_SB_SB1_n643), .A4(R2_SB_SB1_n642), .ZN(R2_SB_n333) );
  NAND3_X1 R2_SB_SB1_U437 ( .A1(R2_SB_SB1_n684), .A2(R2_SB_SB1_n843), .A3(
        R2_SB_SB1_n744), .ZN(R2_SB_SB1_n660) );
  NAND3_X1 R2_SB_SB1_U436 ( .A1(R2_SB_n337), .A2(R2_SB_SB1_n854), .A3(
        R2_SB_SB1_n792), .ZN(R2_SB_SB1_n658) );
  NAND4_X1 R2_SB_SB1_U435 ( .A1(R2_SB_SB1_n660), .A2(R2_SB_SB1_n659), .A3(
        R2_SB_SB1_n658), .A4(R2_SB_SB1_n657), .ZN(R2_SB_SB1_n668) );
  OAI33_X1 R2_SB_SB1_U434 ( .A1(R2_SB_SB1_n862), .A2(R2_SB_n344), .A3(
        R2_SB_SB1_n847), .B1(R2_SB_SB1_n903), .B2(R2_SB_SB1_n858), .B3(
        R2_SB_SB1_n830), .ZN(R2_SB_SB1_n661) );
  NAND3_X1 R2_SB_SB1_U433 ( .A1(R2_SB_SB1_n670), .A2(R2_SB_SB1_n669), .A3(
        R2_SB_SB1_n766), .ZN(R2_SB_SB1_n717) );
  NAND4_X1 R2_SB_SB1_U432 ( .A1(R2_SB_SB1_n717), .A2(R2_SB_SB1_n716), .A3(
        R2_SB_SB1_n677), .A4(R2_SB_SB1_n676), .ZN(R2_SB_SB1_n689) );
  OAI33_X1 R2_SB_SB1_U431 ( .A1(R2_SB_SB1_n839), .A2(R2_SB_SB1_n870), .A3(
        R2_SB_SB1_n883), .B1(R2_SB_SB1_n827), .B2(R2_SB_SB1_n685), .B3(
        R2_SB_SB1_n903), .ZN(R2_SB_SB1_n686) );
  NAND4_X1 R2_SB_SB1_U430 ( .A1(R2_SB_SB1_n693), .A2(R2_SB_SB1_n692), .A3(
        R2_SB_SB1_n691), .A4(R2_SB_SB1_n690), .ZN(R2_SB_n334) );
  NAND3_X1 R2_SB_SB1_U429 ( .A1(R2_SB_SB1_n845), .A2(R2_SB_SB1_n838), .A3(
        R2_SB_SB1_n829), .ZN(R2_SB_SB1_n703) );
  OAI33_X1 R2_SB_SB1_U428 ( .A1(R2_SB_SB1_n876), .A2(R2_SB_n337), .A3(
        R2_SB_SB1_n830), .B1(R2_SB_SB1_n705), .B2(R2_SB_SB1_n835), .B3(
        R2_SB_SB1_n901), .ZN(R2_SB_SB1_n706) );
  NAND3_X1 R2_SB_SB1_U427 ( .A1(R2_SB_n341), .A2(R2_SB_SB1_n714), .A3(
        R2_SB_n344), .ZN(R2_SB_SB1_n715) );
  NAND3_X1 R2_SB_SB1_U426 ( .A1(R2_SB_SB1_n717), .A2(R2_SB_SB1_n716), .A3(
        R2_SB_SB1_n715), .ZN(R2_SB_SB1_n737) );
  NAND4_X1 R2_SB_SB1_U425 ( .A1(R2_SB_SB1_n741), .A2(R2_SB_SB1_n740), .A3(
        R2_SB_SB1_n739), .A4(R2_SB_SB1_n738), .ZN(R2_SB_n335) );
  NAND3_X1 R2_SB_SB1_U424 ( .A1(R2_SB_n344), .A2(R2_SB_SB1_n854), .A3(
        R2_SB_SB1_n795), .ZN(R2_SB_SB1_n762) );
  NAND3_X1 R2_SB_SB1_U423 ( .A1(R2_SB_SB1_n763), .A2(R2_SB_SB1_n762), .A3(
        R2_SB_SB1_n761), .ZN(R2_SB_SB1_n764) );
  NAND3_X1 R2_SB_SB1_U422 ( .A1(R2_SB_n343), .A2(R2_SB_SB1_n854), .A3(
        R2_SB_SB1_n771), .ZN(R2_SB_SB1_n777) );
  NAND3_X1 R2_SB_SB1_U421 ( .A1(R2_SB_SB1_n817), .A2(R2_SB_SB1_n816), .A3(
        R2_SB_SB1_n815), .ZN(R2_SB_SB1_n820) );
  NAND4_X1 R2_SB_SB1_U420 ( .A1(R2_SB_SB1_n825), .A2(R2_SB_SB1_n824), .A3(
        R2_SB_SB1_n823), .A4(R2_SB_SB1_n822), .ZN(R2_SB_n336) );
  NOR2_X2 R2_SB_SB1_U264 ( .A1(R2_SB_SB1_n830), .A2(R2_SB_SB1_n843), .ZN(
        R2_SB_SB1_n758) );
  INV_X1 R2_SB_SB2_U466 ( .A(R2_SB_SB2_n453), .ZN(R2_SB_SB2_n452) );
  INV_X1 R2_SB_SB2_U465 ( .A(R2_SB_n322), .ZN(R2_SB_SB2_n89) );
  INV_X1 R2_SB_SB2_U419 ( .A(R2_SB_n321), .ZN(R2_SB_SB2_n453) );
  NAND2_X1 R2_SB_SB2_U418 ( .A1(R2_SB_n322), .A2(R2_SB_n327), .ZN(
        R2_SB_SB2_n705) );
  AOI22_X1 R2_SB_SB2_U417 ( .A1(R2_SB_SB2_n779), .A2(R2_SB_SB2_n760), .B1(
        R2_SB_SB2_n877), .B2(R2_SB_SB2_n792), .ZN(R2_SB_SB2_n761) );
  OAI21_X1 R2_SB_SB2_U416 ( .B1(R2_SB_SB2_n759), .B2(R2_SB_SB2_n900), .A(
        R2_SB_SB2_n758), .ZN(R2_SB_SB2_n763) );
  AOI222_X1 R2_SB_SB2_U415 ( .A1(R2_SB_SB2_n742), .A2(R2_SB_n326), .B1(
        R2_SB_SB2_n778), .B2(R2_SB_SB2_n748), .C1(R2_SB_SB2_n747), .C2(
        R2_SB_SB2_n656), .ZN(R2_SB_SB2_n657) );
  NAND2_X1 R2_SB_SB2_U414 ( .A1(R2_SB_SB2_n743), .A2(R2_SB_n328), .ZN(
        R2_SB_SB2_n472) );
  AOI21_X1 R2_SB_SB2_U413 ( .B1(R2_SB_SB2_n835), .B2(R2_SB_SB2_n837), .A(
        R2_SB_SB2_n859), .ZN(R2_SB_SB2_n474) );
  OAI21_X1 R2_SB_SB2_U412 ( .B1(R2_SB_SB2_n474), .B2(R2_SB_SB2_n473), .A(
        R2_SB_SB2_n813), .ZN(R2_SB_SB2_n475) );
  OAI22_X1 R2_SB_SB2_U411 ( .A1(R2_SB_SB2_n829), .A2(R2_SB_SB2_n847), .B1(
        R2_SB_SB2_n845), .B2(R2_SB_SB2_n826), .ZN(R2_SB_SB2_n714) );
  NOR2_X1 R2_SB_SB2_U410 ( .A1(R2_SB_n328), .A2(R2_SB_SB2_n863), .ZN(
        R2_SB_SB2_n535) );
  OAI21_X1 R2_SB_SB2_U409 ( .B1(R2_SB_SB2_n855), .B2(R2_SB_SB2_n829), .A(
        R2_SB_SB2_n745), .ZN(R2_SB_SB2_n746) );
  AOI221_X1 R2_SB_SB2_U408 ( .B1(R2_SB_SB2_n805), .B2(R2_SB_SB2_n748), .C1(
        R2_SB_SB2_n747), .C2(R2_SB_SB2_n780), .A(R2_SB_SB2_n746), .ZN(
        R2_SB_SB2_n749) );
  AOI22_X1 R2_SB_SB2_U407 ( .A1(R2_SB_SB2_n742), .A2(R2_SB_n326), .B1(
        R2_SB_SB2_n778), .B2(R2_SB_SB2_n771), .ZN(R2_SB_SB2_n750) );
  OAI211_X1 R2_SB_SB2_U406 ( .C1(R2_SB_SB2_n828), .C2(R2_SB_SB2_n847), .A(
        R2_SB_SB2_n750), .B(R2_SB_SB2_n749), .ZN(R2_SB_SB2_n751) );
  NOR2_X1 R2_SB_SB2_U405 ( .A1(R2_SB_n326), .A2(R2_SB_SB2_n830), .ZN(
        R2_SB_SB2_n724) );
  NOR2_X1 R2_SB_SB2_U404 ( .A1(R2_SB_SB2_n826), .A2(R2_SB_n324), .ZN(
        R2_SB_SB2_n463) );
  OAI22_X1 R2_SB_SB2_U403 ( .A1(R2_SB_n328), .A2(R2_SB_SB2_n876), .B1(
        R2_SB_SB2_n858), .B2(R2_SB_SB2_n901), .ZN(R2_SB_SB2_n760) );
  NOR3_X1 R2_SB_SB2_U402 ( .A1(R2_SB_SB2_n890), .A2(R2_SB_n326), .A3(
        R2_SB_n322), .ZN(R2_SB_SB2_n613) );
  OAI22_X1 R2_SB_SB2_U401 ( .A1(R2_SB_SB2_n89), .A2(R2_SB_SB2_n898), .B1(
        R2_SB_SB2_n628), .B2(R2_SB_SB2_n907), .ZN(R2_SB_SB2_n614) );
  NOR3_X1 R2_SB_SB2_U400 ( .A1(R2_SB_SB2_n614), .A2(R2_SB_SB2_n722), .A3(
        R2_SB_SB2_n613), .ZN(R2_SB_SB2_n623) );
  NOR3_X1 R2_SB_SB2_U399 ( .A1(R2_SB_SB2_n863), .A2(R2_SB_n328), .A3(
        R2_SB_SB2_n814), .ZN(R2_SB_SB2_n797) );
  AOI22_X1 R2_SB_SB2_U398 ( .A1(R2_SB_SB2_n628), .A2(R2_SB_SB2_n627), .B1(
        R2_SB_n323), .B2(R2_SB_SB2_n730), .ZN(R2_SB_SB2_n630) );
  OAI222_X1 R2_SB_SB2_U397 ( .A1(R2_SB_SB2_n837), .A2(R2_SB_SB2_n573), .B1(
        R2_SB_n321), .B2(R2_SB_SB2_n468), .C1(R2_SB_n322), .C2(R2_SB_SB2_n677), 
        .ZN(R2_SB_SB2_n483) );
  OAI221_X1 R2_SB_SB2_U396 ( .B1(R2_SB_n324), .B2(R2_SB_SB2_n581), .C1(
        R2_SB_SB2_n476), .C2(R2_SB_SB2_n878), .A(R2_SB_SB2_n475), .ZN(
        R2_SB_SB2_n482) );
  OAI22_X1 R2_SB_SB2_U395 ( .A1(R2_SB_SB2_n840), .A2(R2_SB_SB2_n800), .B1(
        R2_SB_SB2_n480), .B2(R2_SB_SB2_n453), .ZN(R2_SB_SB2_n481) );
  NOR4_X1 R2_SB_SB2_U394 ( .A1(R2_SB_SB2_n484), .A2(R2_SB_SB2_n483), .A3(
        R2_SB_SB2_n482), .A4(R2_SB_SB2_n481), .ZN(R2_SB_SB2_n485) );
  NOR2_X1 R2_SB_SB2_U393 ( .A1(R2_SB_SB2_n868), .A2(R2_SB_n328), .ZN(
        R2_SB_SB2_n680) );
  NOR2_X1 R2_SB_SB2_U392 ( .A1(R2_SB_n323), .A2(R2_SB_n325), .ZN(
        R2_SB_SB2_n646) );
  NAND2_X1 R2_SB_SB2_U391 ( .A1(R2_SB_n326), .A2(R2_SB_SB2_n872), .ZN(
        R2_SB_SB2_n770) );
  NOR2_X1 R2_SB_SB2_U390 ( .A1(R2_SB_SB2_n895), .A2(R2_SB_n324), .ZN(
        R2_SB_SB2_n783) );
  NOR2_X1 R2_SB_SB2_U389 ( .A1(R2_SB_n325), .A2(R2_SB_n326), .ZN(
        R2_SB_SB2_n617) );
  NOR2_X1 R2_SB_SB2_U388 ( .A1(R2_SB_SB2_n854), .A2(R2_SB_n323), .ZN(
        R2_SB_SB2_n811) );
  INV_X1 R2_SB_SB2_U387 ( .A(R2_SB_n328), .ZN(R2_SB_SB2_n881) );
  AOI22_X1 R2_SB_SB2_U386 ( .A1(R2_SB_n323), .A2(R2_SB_SB2_n638), .B1(
        R2_SB_SB2_n795), .B2(R2_SB_SB2_n713), .ZN(R2_SB_SB2_n711) );
  NOR2_X1 R2_SB_SB2_U385 ( .A1(R2_SB_SB2_n854), .A2(R2_SB_n326), .ZN(
        R2_SB_SB2_n694) );
  NAND2_X1 R2_SB_SB2_U384 ( .A1(R2_SB_n323), .A2(R2_SB_n326), .ZN(
        R2_SB_SB2_n608) );
  OAI221_X1 R2_SB_SB2_U383 ( .B1(R2_SB_n323), .B2(R2_SB_SB2_n551), .C1(
        R2_SB_SB2_n550), .C2(R2_SB_SB2_n910), .A(R2_SB_SB2_n902), .ZN(
        R2_SB_SB2_n552) );
  OAI221_X1 R2_SB_SB2_U382 ( .B1(R2_SB_SB2_n864), .B2(R2_SB_SB2_n838), .C1(
        R2_SB_SB2_n827), .C2(R2_SB_SB2_n849), .A(R2_SB_SB2_n615), .ZN(
        R2_SB_SB2_n553) );
  OAI221_X1 R2_SB_SB2_U381 ( .B1(R2_SB_SB2_n864), .B2(R2_SB_SB2_n835), .C1(
        R2_SB_SB2_n832), .C2(R2_SB_SB2_n853), .A(R2_SB_SB2_n546), .ZN(
        R2_SB_SB2_n554) );
  AOI221_X1 R2_SB_SB2_U380 ( .B1(R2_SB_SB2_n752), .B2(R2_SB_SB2_n554), .C1(
        R2_SB_SB2_n702), .C2(R2_SB_SB2_n553), .A(R2_SB_SB2_n552), .ZN(
        R2_SB_SB2_n559) );
  OAI22_X1 R2_SB_SB2_U379 ( .A1(R2_SB_SB2_n583), .A2(R2_SB_SB2_n826), .B1(
        R2_SB_SB2_n838), .B2(R2_SB_SB2_n891), .ZN(R2_SB_SB2_n584) );
  OAI211_X1 R2_SB_SB2_U378 ( .C1(R2_SB_SB2_n453), .C2(R2_SB_SB2_n844), .A(
        R2_SB_SB2_n835), .B(R2_SB_SB2_n847), .ZN(R2_SB_SB2_n585) );
  OAI211_X1 R2_SB_SB2_U377 ( .C1(R2_SB_n321), .C2(R2_SB_SB2_n898), .A(
        R2_SB_SB2_n582), .B(R2_SB_SB2_n581), .ZN(R2_SB_SB2_n586) );
  AOI221_X1 R2_SB_SB2_U376 ( .B1(R2_SB_n323), .B2(R2_SB_SB2_n586), .C1(
        R2_SB_SB2_n755), .C2(R2_SB_SB2_n585), .A(R2_SB_SB2_n584), .ZN(
        R2_SB_SB2_n599) );
  OAI221_X1 R2_SB_SB2_U375 ( .B1(R2_SB_SB2_n840), .B2(R2_SB_SB2_n859), .C1(
        R2_SB_SB2_n863), .C2(R2_SB_SB2_n834), .A(R2_SB_SB2_n574), .ZN(
        R2_SB_SB2_n580) );
  OAI22_X1 R2_SB_SB2_U374 ( .A1(R2_SB_n324), .A2(R2_SB_SB2_n578), .B1(
        R2_SB_SB2_n577), .B2(R2_SB_SB2_n831), .ZN(R2_SB_SB2_n579) );
  INV_X1 R2_SB_SB2_U373 ( .A(R2_SB_SB2_n573), .ZN(R2_SB_SB2_n889) );
  AOI221_X1 R2_SB_SB2_U372 ( .B1(R2_SB_SB2_n889), .B2(R2_SB_SB2_n696), .C1(
        R2_SB_SB2_n752), .C2(R2_SB_SB2_n580), .A(R2_SB_SB2_n579), .ZN(
        R2_SB_SB2_n600) );
  NOR2_X1 R2_SB_SB2_U371 ( .A1(R2_SB_n324), .A2(R2_SB_n325), .ZN(
        R2_SB_SB2_n656) );
  INV_X1 R2_SB_SB2_U370 ( .A(R2_SB_n327), .ZN(R2_SB_SB2_n872) );
  NOR3_X1 R2_SB_SB2_U369 ( .A1(R2_SB_SB2_n850), .A2(R2_SB_n325), .A3(
        R2_SB_SB2_n881), .ZN(R2_SB_SB2_n556) );
  NOR2_X1 R2_SB_SB2_U368 ( .A1(R2_SB_SB2_n830), .A2(R2_SB_n325), .ZN(
        R2_SB_SB2_n678) );
  AOI221_X1 R2_SB_SB2_U367 ( .B1(R2_SB_SB2_n806), .B2(R2_SB_SB2_n89), .C1(
        R2_SB_SB2_n805), .C2(R2_SB_SB2_n804), .A(R2_SB_SB2_n803), .ZN(
        R2_SB_SB2_n807) );
  AOI211_X1 R2_SB_SB2_U366 ( .C1(R2_SB_SB2_n799), .C2(R2_SB_SB2_n798), .A(
        R2_SB_SB2_n797), .B(R2_SB_SB2_n796), .ZN(R2_SB_SB2_n808) );
  AOI22_X1 R2_SB_SB2_U365 ( .A1(R2_SB_SB2_n793), .A2(R2_SB_SB2_n792), .B1(
        R2_SB_SB2_n791), .B2(R2_SB_SB2_n790), .ZN(R2_SB_SB2_n809) );
  OAI221_X1 R2_SB_SB2_U364 ( .B1(R2_SB_n327), .B2(R2_SB_SB2_n809), .C1(
        R2_SB_SB2_n808), .C2(R2_SB_SB2_n859), .A(R2_SB_SB2_n807), .ZN(
        R2_SB_SB2_n821) );
  NOR2_X1 R2_SB_SB2_U363 ( .A1(R2_SB_n328), .A2(R2_SB_n325), .ZN(
        R2_SB_SB2_n489) );
  OAI21_X1 R2_SB_SB2_U362 ( .B1(R2_SB_SB2_n864), .B2(R2_SB_SB2_n878), .A(
        R2_SB_SB2_n894), .ZN(R2_SB_SB2_n490) );
  AOI221_X1 R2_SB_SB2_U361 ( .B1(R2_SB_SB2_n779), .B2(R2_SB_SB2_n490), .C1(
        R2_SB_SB2_n489), .C2(R2_SB_SB2_n782), .A(R2_SB_SB2_n756), .ZN(
        R2_SB_SB2_n491) );
  AOI222_X1 R2_SB_SB2_U360 ( .A1(R2_SB_SB2_n789), .A2(R2_SB_SB2_n772), .B1(
        R2_SB_SB2_n646), .B2(R2_SB_SB2_n813), .C1(R2_SB_SB2_n709), .C2(
        R2_SB_SB2_n811), .ZN(R2_SB_SB2_n647) );
  OAI221_X1 R2_SB_SB2_U359 ( .B1(R2_SB_n322), .B2(R2_SB_SB2_n884), .C1(
        R2_SB_SB2_n453), .C2(R2_SB_SB2_n880), .A(R2_SB_SB2_n649), .ZN(
        R2_SB_SB2_n650) );
  OAI221_X1 R2_SB_SB2_U358 ( .B1(R2_SB_n324), .B2(R2_SB_SB2_n648), .C1(
        R2_SB_SB2_n845), .C2(R2_SB_SB2_n868), .A(R2_SB_SB2_n647), .ZN(
        R2_SB_SB2_n652) );
  AOI222_X1 R2_SB_SB2_U357 ( .A1(R2_SB_SB2_n781), .A2(R2_SB_SB2_n652), .B1(
        R2_SB_SB2_n651), .B2(R2_SB_SB2_n730), .C1(R2_SB_SB2_n782), .C2(
        R2_SB_SB2_n650), .ZN(R2_SB_SB2_n693) );
  NOR2_X1 R2_SB_SB2_U356 ( .A1(R2_SB_SB2_n863), .A2(R2_SB_n324), .ZN(
        R2_SB_SB2_n618) );
  NOR3_X1 R2_SB_SB2_U355 ( .A1(R2_SB_SB2_n840), .A2(R2_SB_n327), .A3(
        R2_SB_SB2_n869), .ZN(R2_SB_SB2_n575) );
  AOI221_X1 R2_SB_SB2_U354 ( .B1(R2_SB_SB2_n591), .B2(R2_SB_SB2_n453), .C1(
        R2_SB_SB2_n576), .C2(R2_SB_SB2_n684), .A(R2_SB_SB2_n575), .ZN(
        R2_SB_SB2_n578) );
  OAI211_X1 R2_SB_SB2_U353 ( .C1(R2_SB_n326), .C2(R2_SB_SB2_n848), .A(
        R2_SB_SB2_n860), .B(R2_SB_SB2_n853), .ZN(R2_SB_SB2_n662) );
  OAI21_X1 R2_SB_SB2_U352 ( .B1(R2_SB_SB2_n876), .B2(R2_SB_SB2_n853), .A(
        R2_SB_SB2_n908), .ZN(R2_SB_SB2_n663) );
  AOI221_X1 R2_SB_SB2_U351 ( .B1(R2_SB_SB2_n779), .B2(R2_SB_SB2_n663), .C1(
        R2_SB_SB2_n702), .C2(R2_SB_SB2_n662), .A(R2_SB_SB2_n661), .ZN(
        R2_SB_SB2_n664) );
  OAI222_X1 R2_SB_SB2_U350 ( .A1(R2_SB_SB2_n718), .A2(R2_SB_SB2_n907), .B1(
        R2_SB_SB2_n452), .B2(R2_SB_SB2_n664), .C1(R2_SB_SB2_n832), .C2(
        R2_SB_SB2_n802), .ZN(R2_SB_SB2_n667) );
  NOR3_X1 R2_SB_SB2_U349 ( .A1(R2_SB_SB2_n849), .A2(R2_SB_n328), .A3(
        R2_SB_SB2_n854), .ZN(R2_SB_SB2_n605) );
  OAI22_X1 R2_SB_SB2_U348 ( .A1(R2_SB_n327), .A2(R2_SB_n325), .B1(R2_SB_n326), 
        .B2(R2_SB_SB2_n883), .ZN(R2_SB_SB2_n606) );
  AOI221_X1 R2_SB_SB2_U347 ( .B1(R2_SB_SB2_n755), .B2(R2_SB_SB2_n791), .C1(
        R2_SB_SB2_n758), .C2(R2_SB_SB2_n606), .A(R2_SB_SB2_n605), .ZN(
        R2_SB_SB2_n607) );
  NOR2_X1 R2_SB_SB2_U346 ( .A1(R2_SB_SB2_n452), .A2(R2_SB_n323), .ZN(
        R2_SB_SB2_n794) );
  NOR2_X1 R2_SB_SB2_U345 ( .A1(R2_SB_n326), .A2(R2_SB_n328), .ZN(
        R2_SB_SB2_n709) );
  NOR2_X1 R2_SB_SB2_U344 ( .A1(R2_SB_SB2_n830), .A2(R2_SB_n324), .ZN(
        R2_SB_SB2_n782) );
  NOR3_X1 R2_SB_SB2_U343 ( .A1(R2_SB_SB2_n901), .A2(R2_SB_n327), .A3(
        R2_SB_SB2_n843), .ZN(R2_SB_SB2_n729) );
  AOI221_X1 R2_SB_SB2_U342 ( .B1(R2_SB_SB2_n805), .B2(R2_SB_SB2_n813), .C1(
        R2_SB_SB2_n789), .C2(R2_SB_SB2_n728), .A(R2_SB_SB2_n727), .ZN(
        R2_SB_SB2_n732) );
  AOI211_X1 R2_SB_SB2_U341 ( .C1(R2_SB_SB2_n752), .C2(R2_SB_SB2_n730), .A(
        R2_SB_SB2_n759), .B(R2_SB_SB2_n729), .ZN(R2_SB_SB2_n731) );
  OAI222_X1 R2_SB_SB2_U340 ( .A1(R2_SB_SB2_n733), .A2(R2_SB_SB2_n839), .B1(
        R2_SB_SB2_n732), .B2(R2_SB_SB2_n837), .C1(R2_SB_SB2_n731), .C2(
        R2_SB_SB2_n835), .ZN(R2_SB_SB2_n734) );
  NOR2_X1 R2_SB_SB2_U339 ( .A1(R2_SB_SB2_n854), .A2(R2_SB_n324), .ZN(
        R2_SB_SB2_n805) );
  NOR2_X1 R2_SB_SB2_U338 ( .A1(R2_SB_SB2_n872), .A2(R2_SB_n326), .ZN(
        R2_SB_SB2_n767) );
  INV_X1 R2_SB_SB2_U337 ( .A(R2_SB_n323), .ZN(R2_SB_SB2_n830) );
  NOR2_X1 R2_SB_SB2_U336 ( .A1(R2_SB_n327), .A2(R2_SB_n328), .ZN(
        R2_SB_SB2_n702) );
  NOR2_X1 R2_SB_SB2_U335 ( .A1(R2_SB_n322), .A2(R2_SB_n323), .ZN(
        R2_SB_SB2_n795) );
  NOR2_X1 R2_SB_SB2_U334 ( .A1(R2_SB_n326), .A2(R2_SB_n327), .ZN(
        R2_SB_SB2_n813) );
  NOR3_X1 R2_SB_SB2_U333 ( .A1(R2_SB_SB2_n833), .A2(R2_SB_n324), .A3(
        R2_SB_SB2_n885), .ZN(R2_SB_SB2_n639) );
  INV_X1 R2_SB_SB2_U332 ( .A(R2_SB_n325), .ZN(R2_SB_SB2_n854) );
  NOR2_X1 R2_SB_SB2_U331 ( .A1(R2_SB_SB2_n843), .A2(R2_SB_n323), .ZN(
        R2_SB_SB2_n792) );
  INV_X1 R2_SB_SB2_U330 ( .A(R2_SB_n326), .ZN(R2_SB_SB2_n863) );
  NAND2_X1 R2_SB_SB2_U329 ( .A1(R2_SB_SB2_n791), .A2(R2_SB_SB2_n772), .ZN(
        R2_SB_SB2_n775) );
  OAI21_X1 R2_SB_SB2_U328 ( .B1(R2_SB_SB2_n775), .B2(R2_SB_SB2_n774), .A(
        R2_SB_SB2_n773), .ZN(R2_SB_SB2_n776) );
  INV_X1 R2_SB_SB2_U327 ( .A(R2_SB_SB2_n776), .ZN(R2_SB_SB2_n887) );
  INV_X1 R2_SB_SB2_U326 ( .A(R2_SB_SB2_n783), .ZN(R2_SB_SB2_n897) );
  INV_X1 R2_SB_SB2_U325 ( .A(R2_SB_SB2_n678), .ZN(R2_SB_SB2_n860) );
  INV_X1 R2_SB_SB2_U324 ( .A(R2_SB_SB2_n811), .ZN(R2_SB_SB2_n855) );
  INV_X1 R2_SB_SB2_U323 ( .A(R2_SB_SB2_n463), .ZN(R2_SB_SB2_n842) );
  INV_X1 R2_SB_SB2_U322 ( .A(R2_SB_SB2_n711), .ZN(R2_SB_SB2_n909) );
  NAND2_X1 R2_SB_SB2_U321 ( .A1(R2_SB_SB2_n678), .A2(R2_SB_SB2_n781), .ZN(
        R2_SB_SB2_n615) );
  NAND2_X1 R2_SB_SB2_U320 ( .A1(R2_SB_SB2_n680), .A2(R2_SB_SB2_n810), .ZN(
        R2_SB_SB2_n581) );
  NAND2_X1 R2_SB_SB2_U319 ( .A1(R2_SB_SB2_n772), .A2(R2_SB_SB2_n684), .ZN(
        R2_SB_SB2_n785) );
  NAND2_X1 R2_SB_SB2_U318 ( .A1(R2_SB_SB2_n670), .A2(R2_SB_SB2_n881), .ZN(
        R2_SB_SB2_n773) );
  NAND2_X1 R2_SB_SB2_U317 ( .A1(R2_SB_SB2_n670), .A2(R2_SB_SB2_n872), .ZN(
        R2_SB_SB2_n801) );
  NAND2_X1 R2_SB_SB2_U316 ( .A1(R2_SB_SB2_n452), .A2(R2_SB_SB2_n843), .ZN(
        R2_SB_SB2_n548) );
  NOR2_X1 R2_SB_SB2_U315 ( .A1(R2_SB_SB2_n854), .A2(R2_SB_SB2_n827), .ZN(
        R2_SB_SB2_n793) );
  OAI21_X1 R2_SB_SB2_U314 ( .B1(R2_SB_SB2_n718), .B2(R2_SB_SB2_n588), .A(
        R2_SB_SB2_n587), .ZN(R2_SB_SB2_n597) );
  AOI22_X1 R2_SB_SB2_U313 ( .A1(R2_SB_SB2_n753), .A2(R2_SB_SB2_n771), .B1(
        R2_SB_SB2_n752), .B2(R2_SB_SB2_n751), .ZN(R2_SB_SB2_n825) );
  AOI22_X1 R2_SB_SB2_U312 ( .A1(R2_SB_n322), .A2(R2_SB_SB2_n765), .B1(
        R2_SB_SB2_n764), .B2(R2_SB_SB2_n453), .ZN(R2_SB_SB2_n824) );
  NOR4_X1 R2_SB_SB2_U311 ( .A1(R2_SB_SB2_n464), .A2(R2_SB_SB2_n886), .A3(
        R2_SB_SB2_n555), .A4(R2_SB_SB2_n639), .ZN(R2_SB_SB2_n486) );
  AOI211_X1 R2_SB_SB2_U310 ( .C1(R2_SB_SB2_n684), .C2(R2_SB_SB2_n462), .A(
        R2_SB_SB2_n461), .B(R2_SB_SB2_n460), .ZN(R2_SB_SB2_n487) );
  AOI221_X1 R2_SB_SB2_U309 ( .B1(R2_SB_SB2_n810), .B2(R2_SB_SB2_n533), .C1(
        R2_SB_SB2_n565), .C2(R2_SB_n322), .A(R2_SB_SB2_n532), .ZN(
        R2_SB_SB2_n561) );
  NOR4_X1 R2_SB_SB2_U308 ( .A1(R2_SB_SB2_n557), .A2(R2_SB_SB2_n556), .A3(
        R2_SB_SB2_n555), .A4(R2_SB_SB2_n674), .ZN(R2_SB_SB2_n558) );
  AOI221_X1 R2_SB_SB2_U307 ( .B1(R2_SB_SB2_n772), .B2(R2_SB_SB2_n572), .C1(
        R2_SB_SB2_n753), .C2(R2_SB_SB2_n758), .A(R2_SB_SB2_n571), .ZN(
        R2_SB_SB2_n601) );
  AOI211_X1 R2_SB_SB2_U306 ( .C1(R2_SB_SB2_n597), .C2(R2_SB_SB2_n453), .A(
        R2_SB_SB2_n596), .B(R2_SB_SB2_n595), .ZN(R2_SB_SB2_n598) );
  AOI221_X1 R2_SB_SB2_U305 ( .B1(R2_SB_SB2_n604), .B2(R2_SB_SB2_n877), .C1(
        R2_SB_SB2_n603), .C2(R2_SB_SB2_n679), .A(R2_SB_SB2_n602), .ZN(
        R2_SB_SB2_n645) );
  NOR4_X1 R2_SB_SB2_U304 ( .A1(R2_SB_SB2_n641), .A2(R2_SB_SB2_n640), .A3(
        R2_SB_SB2_n639), .A4(R2_SB_SB2_n673), .ZN(R2_SB_SB2_n642) );
  OAI21_X1 R2_SB_SB2_U303 ( .B1(R2_SB_SB2_n810), .B2(R2_SB_SB2_n744), .A(
        R2_SB_SB2_n743), .ZN(R2_SB_SB2_n745) );
  NOR4_X1 R2_SB_SB2_U302 ( .A1(R2_SB_SB2_n737), .A2(R2_SB_SB2_n736), .A3(
        R2_SB_SB2_n735), .A4(R2_SB_SB2_n734), .ZN(R2_SB_SB2_n738) );
  AOI211_X1 R2_SB_SB2_U301 ( .C1(R2_SB_SB2_n713), .C2(R2_SB_SB2_n758), .A(
        R2_SB_SB2_n712), .B(R2_SB_SB2_n909), .ZN(R2_SB_SB2_n739) );
  NOR4_X1 R2_SB_SB2_U300 ( .A1(R2_SB_SB2_n689), .A2(R2_SB_SB2_n688), .A3(
        R2_SB_SB2_n687), .A4(R2_SB_SB2_n686), .ZN(R2_SB_SB2_n690) );
  AOI211_X1 R2_SB_SB2_U299 ( .C1(R2_SB_SB2_n752), .C2(R2_SB_SB2_n668), .A(
        R2_SB_SB2_n667), .B(R2_SB_SB2_n666), .ZN(R2_SB_SB2_n691) );
  AOI221_X1 R2_SB_SB2_U298 ( .B1(R2_SB_SB2_n565), .B2(R2_SB_SB2_n766), .C1(
        R2_SB_SB2_n759), .C2(R2_SB_SB2_n791), .A(R2_SB_SB2_n513), .ZN(
        R2_SB_SB2_n525) );
  NOR4_X1 R2_SB_SB2_U297 ( .A1(R2_SB_SB2_n523), .A2(R2_SB_SB2_n522), .A3(
        R2_SB_SB2_n521), .A4(R2_SB_SB2_n520), .ZN(R2_SB_SB2_n524) );
  OAI221_X1 R2_SB_SB2_U296 ( .B1(R2_SB_SB2_n849), .B2(R2_SB_SB2_n770), .C1(
        R2_SB_SB2_n883), .C2(R2_SB_SB2_n608), .A(R2_SB_SB2_n567), .ZN(
        R2_SB_SB2_n568) );
  OAI21_X1 R2_SB_SB2_U295 ( .B1(R2_SB_SB2_n569), .B2(R2_SB_SB2_n568), .A(
        R2_SB_SB2_n781), .ZN(R2_SB_SB2_n570) );
  OAI21_X1 R2_SB_SB2_U294 ( .B1(R2_SB_SB2_n839), .B2(R2_SB_SB2_n892), .A(
        R2_SB_SB2_n570), .ZN(R2_SB_SB2_n571) );
  INV_X1 R2_SB_SB2_U293 ( .A(R2_SB_SB2_n780), .ZN(R2_SB_SB2_n870) );
  OAI21_X1 R2_SB_SB2_U292 ( .B1(R2_SB_SB2_n778), .B2(R2_SB_SB2_n744), .A(
        R2_SB_SB2_n696), .ZN(R2_SB_SB2_n508) );
  OAI211_X1 R2_SB_SB2_U291 ( .C1(R2_SB_SB2_n813), .C2(R2_SB_SB2_n812), .A(
        R2_SB_SB2_n811), .B(R2_SB_SB2_n810), .ZN(R2_SB_SB2_n817) );
  INV_X1 R2_SB_SB2_U290 ( .A(R2_SB_SB2_n743), .ZN(R2_SB_SB2_n851) );
  AND3_X1 R2_SB_SB2_U289 ( .A1(R2_SB_SB2_n779), .A2(R2_SB_SB2_n812), .A3(
        R2_SB_SB2_n656), .ZN(R2_SB_SB2_n87) );
  NOR3_X1 R2_SB_SB2_U288 ( .A1(R2_SB_SB2_n858), .A2(R2_SB_SB2_n665), .A3(
        R2_SB_SB2_n890), .ZN(R2_SB_SB2_n13) );
  OR3_X1 R2_SB_SB2_U287 ( .A1(R2_SB_SB2_n13), .A2(R2_SB_SB2_n675), .A3(
        R2_SB_SB2_n87), .ZN(R2_SB_SB2_n464) );
  OAI22_X1 R2_SB_SB2_U286 ( .A1(R2_SB_SB2_n872), .A2(R2_SB_SB2_n857), .B1(
        R2_SB_SB2_n854), .B2(R2_SB_SB2_n876), .ZN(R2_SB_SB2_n547) );
  INV_X1 R2_SB_SB2_U285 ( .A(R2_SB_SB2_n582), .ZN(R2_SB_SB2_n911) );
  AOI21_X1 R2_SB_SB2_U284 ( .B1(R2_SB_SB2_n781), .B2(R2_SB_SB2_n547), .A(
        R2_SB_SB2_n911), .ZN(R2_SB_SB2_n551) );
  AOI21_X1 R2_SB_SB2_U283 ( .B1(R2_SB_SB2_n754), .B2(R2_SB_SB2_n758), .A(
        R2_SB_SB2_n467), .ZN(R2_SB_SB2_n468) );
  AOI21_X1 R2_SB_SB2_U282 ( .B1(R2_SB_SB2_n778), .B2(R2_SB_SB2_n453), .A(
        R2_SB_SB2_n789), .ZN(R2_SB_SB2_n700) );
  AOI22_X1 R2_SB_SB2_U281 ( .A1(R2_SB_SB2_n725), .A2(R2_SB_SB2_n617), .B1(
        R2_SB_SB2_n766), .B2(R2_SB_SB2_n730), .ZN(R2_SB_SB2_n562) );
  AOI21_X1 R2_SB_SB2_U280 ( .B1(R2_SB_SB2_n743), .B2(R2_SB_n322), .A(
        R2_SB_SB2_n747), .ZN(R2_SB_SB2_n564) );
  OAI21_X1 R2_SB_SB2_U279 ( .B1(R2_SB_SB2_n684), .B2(R2_SB_SB2_n799), .A(
        R2_SB_SB2_n780), .ZN(R2_SB_SB2_n563) );
  OAI211_X1 R2_SB_SB2_U278 ( .C1(R2_SB_SB2_n564), .C2(R2_SB_SB2_n868), .A(
        R2_SB_SB2_n563), .B(R2_SB_SB2_n562), .ZN(R2_SB_SB2_n572) );
  OAI21_X1 R2_SB_SB2_U277 ( .B1(R2_SB_SB2_n905), .B2(R2_SB_SB2_n859), .A(
        R2_SB_SB2_n895), .ZN(R2_SB_SB2_n529) );
  AOI211_X1 R2_SB_SB2_U276 ( .C1(R2_SB_SB2_n529), .C2(R2_SB_SB2_n830), .A(
        R2_SB_SB2_n633), .B(R2_SB_SB2_n528), .ZN(R2_SB_SB2_n530) );
  AOI22_X1 R2_SB_SB2_U275 ( .A1(R2_SB_SB2_n680), .A2(R2_SB_SB2_n843), .B1(
        R2_SB_SB2_n678), .B2(R2_SB_SB2_n772), .ZN(R2_SB_SB2_n531) );
  OAI211_X1 R2_SB_SB2_U274 ( .C1(R2_SB_SB2_n905), .C2(R2_SB_SB2_n864), .A(
        R2_SB_SB2_n531), .B(R2_SB_SB2_n530), .ZN(R2_SB_SB2_n533) );
  OAI21_X1 R2_SB_SB2_U273 ( .B1(R2_SB_SB2_n755), .B2(R2_SB_SB2_n754), .A(
        R2_SB_SB2_n782), .ZN(R2_SB_SB2_n757) );
  INV_X1 R2_SB_SB2_U272 ( .A(R2_SB_SB2_n756), .ZN(R2_SB_SB2_n899) );
  OAI211_X1 R2_SB_SB2_U271 ( .C1(R2_SB_SB2_n845), .C2(R2_SB_SB2_n880), .A(
        R2_SB_SB2_n757), .B(R2_SB_SB2_n899), .ZN(R2_SB_SB2_n765) );
  INV_X1 R2_SB_SB2_U270 ( .A(R2_SB_SB2_n696), .ZN(R2_SB_SB2_n836) );
  AOI21_X1 R2_SB_SB2_U269 ( .B1(R2_SB_SB2_n843), .B2(R2_SB_SB2_n835), .A(
        R2_SB_SB2_n879), .ZN(R2_SB_SB2_n595) );
  NAND2_X1 R2_SB_SB2_U268 ( .A1(R2_SB_SB2_n634), .A2(R2_SB_SB2_n805), .ZN(
        R2_SB_SB2_n800) );
  NAND2_X1 R2_SB_SB2_U267 ( .A1(R2_SB_SB2_n772), .A2(R2_SB_SB2_n507), .ZN(
        R2_SB_SB2_n648) );
  AOI21_X1 R2_SB_SB2_U266 ( .B1(R2_SB_SB2_n849), .B2(R2_SB_SB2_n608), .A(
        R2_SB_SB2_n878), .ZN(R2_SB_SB2_n528) );
  INV_X1 R2_SB_SB2_U265 ( .A(R2_SB_SB2_n794), .ZN(R2_SB_SB2_n837) );
  NOR2_X1 R2_SB_SB2_U263 ( .A1(R2_SB_SB2_n770), .A2(R2_SB_SB2_n833), .ZN(
        R2_SB_SB2_n651) );
  INV_X1 R2_SB_SB2_U262 ( .A(R2_SB_SB2_n798), .ZN(R2_SB_SB2_n901) );
  INV_X1 R2_SB_SB2_U261 ( .A(R2_SB_SB2_n813), .ZN(R2_SB_SB2_n876) );
  AOI22_X1 R2_SB_SB2_U260 ( .A1(R2_SB_SB2_n696), .A2(R2_SB_SB2_n789), .B1(
        R2_SB_SB2_n778), .B2(R2_SB_SB2_n779), .ZN(R2_SB_SB2_n612) );
  AOI22_X1 R2_SB_SB2_U259 ( .A1(R2_SB_SB2_n795), .A2(R2_SB_SB2_n798), .B1(
        R2_SB_SB2_n767), .B2(R2_SB_SB2_n766), .ZN(R2_SB_SB2_n768) );
  NAND2_X1 R2_SB_SB2_U258 ( .A1(R2_SB_SB2_n865), .A2(R2_SB_SB2_n853), .ZN(
        R2_SB_SB2_n495) );
  AOI22_X1 R2_SB_SB2_U257 ( .A1(R2_SB_SB2_n684), .A2(R2_SB_SB2_n495), .B1(
        R2_SB_SB2_n696), .B2(R2_SB_SB2_n618), .ZN(R2_SB_SB2_n496) );
  INV_X1 R2_SB_SB2_U256 ( .A(R2_SB_SB2_n805), .ZN(R2_SB_SB2_n857) );
  NAND2_X1 R2_SB_SB2_U255 ( .A1(R2_SB_SB2_n843), .A2(R2_SB_SB2_n863), .ZN(
        R2_SB_SB2_n774) );
  AOI22_X1 R2_SB_SB2_U254 ( .A1(R2_SB_SB2_n798), .A2(R2_SB_SB2_n627), .B1(
        R2_SB_SB2_n743), .B2(R2_SB_SB2_n752), .ZN(R2_SB_SB2_n567) );
  INV_X1 R2_SB_SB2_U253 ( .A(R2_SB_SB2_n767), .ZN(R2_SB_SB2_n874) );
  NOR2_X1 R2_SB_SB2_U252 ( .A1(R2_SB_SB2_n795), .A2(R2_SB_SB2_n794), .ZN(
        R2_SB_SB2_n814) );
  INV_X1 R2_SB_SB2_U251 ( .A(R2_SB_SB2_n694), .ZN(R2_SB_SB2_n869) );
  NOR2_X1 R2_SB_SB2_U250 ( .A1(R2_SB_SB2_n830), .A2(R2_SB_SB2_n684), .ZN(
        R2_SB_SB2_n665) );
  NOR2_X1 R2_SB_SB2_U249 ( .A1(R2_SB_SB2_n843), .A2(R2_SB_n322), .ZN(
        R2_SB_SB2_n604) );
  NOR2_X1 R2_SB_SB2_U248 ( .A1(R2_SB_SB2_n863), .A2(R2_SB_SB2_n858), .ZN(
        R2_SB_SB2_n790) );
  NAND2_X1 R2_SB_SB2_U247 ( .A1(R2_SB_SB2_n752), .A2(R2_SB_SB2_n507), .ZN(
        R2_SB_SB2_n802) );
  AOI21_X1 R2_SB_SB2_U246 ( .B1(R2_SB_SB2_n789), .B2(R2_SB_SB2_n798), .A(
        R2_SB_SB2_n783), .ZN(R2_SB_SB2_n721) );
  OAI21_X1 R2_SB_SB2_U245 ( .B1(R2_SB_SB2_n747), .B2(R2_SB_SB2_n843), .A(
        R2_SB_SB2_n759), .ZN(R2_SB_SB2_n719) );
  OR3_X1 R2_SB_SB2_U244 ( .A1(R2_SB_SB2_n718), .A2(R2_SB_SB2_n452), .A3(
        R2_SB_SB2_n802), .ZN(R2_SB_SB2_n720) );
  OAI211_X1 R2_SB_SB2_U243 ( .C1(R2_SB_SB2_n721), .C2(R2_SB_SB2_n826), .A(
        R2_SB_SB2_n720), .B(R2_SB_SB2_n719), .ZN(R2_SB_SB2_n736) );
  AOI22_X1 R2_SB_SB2_U242 ( .A1(R2_SB_SB2_n678), .A2(R2_SB_SB2_n767), .B1(
        R2_SB_SB2_n900), .B2(R2_SB_SB2_n843), .ZN(R2_SB_SB2_n683) );
  OAI21_X1 R2_SB_SB2_U241 ( .B1(R2_SB_SB2_n794), .B2(R2_SB_SB2_n791), .A(
        R2_SB_SB2_n882), .ZN(R2_SB_SB2_n681) );
  OAI21_X1 R2_SB_SB2_U240 ( .B1(R2_SB_SB2_n680), .B2(R2_SB_SB2_n679), .A(
        R2_SB_SB2_n696), .ZN(R2_SB_SB2_n682) );
  OAI211_X1 R2_SB_SB2_U239 ( .C1(R2_SB_SB2_n683), .C2(R2_SB_SB2_n829), .A(
        R2_SB_SB2_n682), .B(R2_SB_SB2_n681), .ZN(R2_SB_SB2_n688) );
  NOR3_X1 R2_SB_SB2_U238 ( .A1(R2_SB_SB2_n848), .A2(R2_SB_SB2_n452), .A3(
        R2_SB_SB2_n863), .ZN(R2_SB_SB2_n540) );
  OAI22_X1 R2_SB_SB2_U237 ( .A1(R2_SB_SB2_n858), .A2(R2_SB_SB2_n838), .B1(
        R2_SB_SB2_n857), .B2(R2_SB_SB2_n840), .ZN(R2_SB_SB2_n541) );
  AOI21_X1 R2_SB_SB2_U236 ( .B1(R2_SB_n322), .B2(R2_SB_SB2_n548), .A(
        R2_SB_SB2_n862), .ZN(R2_SB_SB2_n539) );
  NOR3_X1 R2_SB_SB2_U235 ( .A1(R2_SB_SB2_n541), .A2(R2_SB_SB2_n540), .A3(
        R2_SB_SB2_n539), .ZN(R2_SB_SB2_n542) );
  AOI21_X1 R2_SB_SB2_U234 ( .B1(R2_SB_SB2_n730), .B2(R2_SB_SB2_n709), .A(
        R2_SB_SB2_n753), .ZN(R2_SB_SB2_n733) );
  INV_X1 R2_SB_SB2_U233 ( .A(R2_SB_SB2_n791), .ZN(R2_SB_SB2_n840) );
  NOR3_X1 R2_SB_SB2_U232 ( .A1(R2_SB_SB2_n828), .A2(R2_SB_SB2_n856), .A3(
        R2_SB_SB2_n876), .ZN(R2_SB_SB2_n819) );
  AOI21_X1 R2_SB_SB2_U231 ( .B1(R2_SB_SB2_n845), .B2(R2_SB_SB2_n837), .A(
        R2_SB_SB2_n906), .ZN(R2_SB_SB2_n818) );
  NOR4_X1 R2_SB_SB2_U230 ( .A1(R2_SB_SB2_n821), .A2(R2_SB_SB2_n820), .A3(
        R2_SB_SB2_n819), .A4(R2_SB_SB2_n818), .ZN(R2_SB_SB2_n822) );
  INV_X1 R2_SB_SB2_U229 ( .A(R2_SB_SB2_n789), .ZN(R2_SB_SB2_n853) );
  NOR2_X1 R2_SB_SB2_U228 ( .A1(R2_SB_SB2_n743), .A2(R2_SB_SB2_n603), .ZN(
        R2_SB_SB2_n718) );
  AOI221_X1 R2_SB_SB2_U227 ( .B1(R2_SB_SB2_n877), .B2(R2_SB_SB2_n684), .C1(
        R2_SB_SB2_n591), .C2(R2_SB_SB2_n89), .A(R2_SB_SB2_n590), .ZN(
        R2_SB_SB2_n593) );
  AOI22_X1 R2_SB_SB2_U226 ( .A1(R2_SB_SB2_n810), .A2(R2_SB_SB2_n589), .B1(
        R2_SB_SB2_n798), .B2(R2_SB_SB2_n723), .ZN(R2_SB_SB2_n594) );
  OAI221_X1 R2_SB_SB2_U225 ( .B1(R2_SB_SB2_n594), .B2(R2_SB_SB2_n859), .C1(
        R2_SB_SB2_n593), .C2(R2_SB_SB2_n849), .A(R2_SB_SB2_n592), .ZN(
        R2_SB_SB2_n596) );
  INV_X1 R2_SB_SB2_U224 ( .A(R2_SB_SB2_n744), .ZN(R2_SB_SB2_n868) );
  OAI21_X1 R2_SB_SB2_U223 ( .B1(R2_SB_SB2_n779), .B2(R2_SB_SB2_n453), .A(
        R2_SB_SB2_n656), .ZN(R2_SB_SB2_n503) );
  NOR2_X1 R2_SB_SB2_U222 ( .A1(R2_SB_SB2_n618), .A2(R2_SB_SB2_n780), .ZN(
        R2_SB_SB2_n504) );
  OAI221_X1 R2_SB_SB2_U221 ( .B1(R2_SB_SB2_n504), .B2(R2_SB_SB2_n840), .C1(
        R2_SB_SB2_n869), .C2(R2_SB_SB2_n852), .A(R2_SB_SB2_n503), .ZN(
        R2_SB_SB2_n505) );
  INV_X1 R2_SB_SB2_U220 ( .A(R2_SB_SB2_n617), .ZN(R2_SB_SB2_n862) );
  AOI21_X1 R2_SB_SB2_U219 ( .B1(R2_SB_SB2_n828), .B2(R2_SB_SB2_n850), .A(
        R2_SB_SB2_n879), .ZN(R2_SB_SB2_n459) );
  AOI221_X1 R2_SB_SB2_U218 ( .B1(R2_SB_SB2_n463), .B2(R2_SB_SB2_n591), .C1(
        R2_SB_SB2_n514), .C2(R2_SB_SB2_n766), .A(R2_SB_SB2_n459), .ZN(
        R2_SB_SB2_n488) );
  OAI222_X1 R2_SB_SB2_U217 ( .A1(R2_SB_SB2_n623), .A2(R2_SB_SB2_n851), .B1(
        R2_SB_SB2_n622), .B2(R2_SB_SB2_n883), .C1(R2_SB_SB2_n621), .C2(
        R2_SB_SB2_n905), .ZN(R2_SB_SB2_n624) );
  OAI221_X1 R2_SB_SB2_U216 ( .B1(R2_SB_SB2_n903), .B2(R2_SB_SB2_n844), .C1(
        R2_SB_SB2_n848), .C2(R2_SB_SB2_n910), .A(R2_SB_SB2_n607), .ZN(
        R2_SB_SB2_n626) );
  OAI211_X1 R2_SB_SB2_U215 ( .C1(R2_SB_SB2_n857), .C2(R2_SB_SB2_n831), .A(
        R2_SB_SB2_n612), .B(R2_SB_SB2_n611), .ZN(R2_SB_SB2_n625) );
  AOI221_X1 R2_SB_SB2_U214 ( .B1(R2_SB_SB2_n452), .B2(R2_SB_SB2_n626), .C1(
        R2_SB_SB2_n752), .C2(R2_SB_SB2_n625), .A(R2_SB_SB2_n624), .ZN(
        R2_SB_SB2_n644) );
  OAI22_X1 R2_SB_SB2_U213 ( .A1(R2_SB_SB2_n733), .A2(R2_SB_SB2_n837), .B1(
        R2_SB_SB2_n842), .B2(R2_SB_SB2_n884), .ZN(R2_SB_SB2_n653) );
  OAI22_X1 R2_SB_SB2_U212 ( .A1(R2_SB_SB2_n858), .A2(R2_SB_SB2_n834), .B1(
        R2_SB_n322), .B2(R2_SB_SB2_n859), .ZN(R2_SB_SB2_n654) );
  OAI21_X1 R2_SB_SB2_U211 ( .B1(R2_SB_SB2_n903), .B2(R2_SB_SB2_n859), .A(
        R2_SB_SB2_n895), .ZN(R2_SB_SB2_n655) );
  AOI221_X1 R2_SB_SB2_U210 ( .B1(R2_SB_SB2_n795), .B2(R2_SB_SB2_n655), .C1(
        R2_SB_SB2_n702), .C2(R2_SB_SB2_n654), .A(R2_SB_SB2_n653), .ZN(
        R2_SB_SB2_n692) );
  AOI221_X1 R2_SB_SB2_U209 ( .B1(R2_SB_SB2_n684), .B2(R2_SB_SB2_n536), .C1(
        R2_SB_SB2_n535), .C2(R2_SB_SB2_n628), .A(R2_SB_SB2_n534), .ZN(
        R2_SB_SB2_n537) );
  OAI222_X1 R2_SB_SB2_U208 ( .A1(R2_SB_SB2_n543), .A2(R2_SB_SB2_n847), .B1(
        R2_SB_SB2_n835), .B2(R2_SB_SB2_n573), .C1(R2_SB_SB2_n542), .C2(
        R2_SB_SB2_n883), .ZN(R2_SB_SB2_n544) );
  OAI221_X1 R2_SB_SB2_U207 ( .B1(R2_SB_SB2_n89), .B2(R2_SB_SB2_n588), .C1(
        R2_SB_n321), .C2(R2_SB_SB2_n910), .A(R2_SB_SB2_n537), .ZN(
        R2_SB_SB2_n545) );
  AOI221_X1 R2_SB_SB2_U206 ( .B1(R2_SB_SB2_n792), .B2(R2_SB_SB2_n545), .C1(
        R2_SB_SB2_n753), .C2(R2_SB_SB2_n791), .A(R2_SB_SB2_n544), .ZN(
        R2_SB_SB2_n560) );
  AOI22_X1 R2_SB_SB2_U205 ( .A1(R2_SB_SB2_n798), .A2(R2_SB_SB2_n708), .B1(
        R2_SB_SB2_n795), .B2(R2_SB_SB2_n767), .ZN(R2_SB_SB2_n631) );
  AOI21_X1 R2_SB_SB2_U204 ( .B1(R2_SB_SB2_n755), .B2(R2_SB_SB2_n758), .A(
        R2_SB_SB2_n756), .ZN(R2_SB_SB2_n629) );
  OAI222_X1 R2_SB_SB2_U203 ( .A1(R2_SB_SB2_n631), .A2(R2_SB_SB2_n857), .B1(
        R2_SB_SB2_n630), .B2(R2_SB_SB2_n875), .C1(R2_SB_n322), .C2(
        R2_SB_SB2_n629), .ZN(R2_SB_SB2_n632) );
  AOI221_X1 R2_SB_SB2_U202 ( .B1(R2_SB_SB2_n725), .B2(R2_SB_SB2_n728), .C1(
        R2_SB_SB2_n651), .C2(R2_SB_SB2_n789), .A(R2_SB_SB2_n632), .ZN(
        R2_SB_SB2_n643) );
  OAI222_X1 R2_SB_SB2_U201 ( .A1(R2_SB_SB2_n865), .A2(R2_SB_SB2_n785), .B1(
        R2_SB_SB2_n784), .B2(R2_SB_SB2_n905), .C1(R2_SB_SB2_n827), .C2(
        R2_SB_SB2_n897), .ZN(R2_SB_SB2_n786) );
  OAI211_X1 R2_SB_SB2_U200 ( .C1(R2_SB_SB2_n829), .C2(R2_SB_SB2_n770), .A(
        R2_SB_SB2_n769), .B(R2_SB_SB2_n768), .ZN(R2_SB_SB2_n788) );
  OAI211_X1 R2_SB_SB2_U199 ( .C1(R2_SB_SB2_n895), .C2(R2_SB_SB2_n848), .A(
        R2_SB_SB2_n777), .B(R2_SB_SB2_n887), .ZN(R2_SB_SB2_n787) );
  AOI221_X1 R2_SB_SB2_U198 ( .B1(R2_SB_SB2_n789), .B2(R2_SB_SB2_n788), .C1(
        R2_SB_n321), .C2(R2_SB_SB2_n787), .A(R2_SB_SB2_n786), .ZN(
        R2_SB_SB2_n823) );
  INV_X1 R2_SB_SB2_U197 ( .A(R2_SB_SB2_n656), .ZN(R2_SB_SB2_n859) );
  AOI211_X1 R2_SB_SB2_U196 ( .C1(R2_SB_SB2_n789), .C2(R2_SB_SB2_n812), .A(
        R2_SB_SB2_n882), .B(R2_SB_SB2_n727), .ZN(R2_SB_SB2_n577) );
  AOI211_X1 R2_SB_SB2_U195 ( .C1(R2_SB_SB2_n744), .C2(R2_SB_SB2_n843), .A(
        R2_SB_SB2_n730), .B(R2_SB_SB2_n792), .ZN(R2_SB_SB2_n509) );
  AOI21_X1 R2_SB_SB2_U194 ( .B1(R2_SB_SB2_n854), .B2(R2_SB_SB2_n881), .A(
        R2_SB_SB2_n767), .ZN(R2_SB_SB2_n477) );
  OAI222_X1 R2_SB_SB2_U193 ( .A1(R2_SB_SB2_n843), .A2(R2_SB_SB2_n885), .B1(
        R2_SB_SB2_n477), .B2(R2_SB_SB2_n845), .C1(R2_SB_SB2_n864), .C2(
        R2_SB_SB2_n878), .ZN(R2_SB_SB2_n479) );
  OAI22_X1 R2_SB_SB2_U192 ( .A1(R2_SB_SB2_n849), .A2(R2_SB_SB2_n648), .B1(
        R2_SB_SB2_n862), .B2(R2_SB_SB2_n844), .ZN(R2_SB_SB2_n478) );
  AOI211_X1 R2_SB_SB2_U191 ( .C1(R2_SB_SB2_n791), .C2(R2_SB_SB2_n812), .A(
        R2_SB_SB2_n479), .B(R2_SB_SB2_n478), .ZN(R2_SB_SB2_n480) );
  NOR3_X1 R2_SB_SB2_U190 ( .A1(R2_SB_SB2_n838), .A2(R2_SB_n321), .A3(
        R2_SB_SB2_n864), .ZN(R2_SB_SB2_n610) );
  AOI21_X1 R2_SB_SB2_U189 ( .B1(R2_SB_SB2_n858), .B2(R2_SB_SB2_n608), .A(
        R2_SB_SB2_n827), .ZN(R2_SB_SB2_n609) );
  AOI211_X1 R2_SB_SB2_U188 ( .C1(R2_SB_SB2_n646), .C2(R2_SB_SB2_n781), .A(
        R2_SB_SB2_n610), .B(R2_SB_SB2_n609), .ZN(R2_SB_SB2_n611) );
  INV_X1 R2_SB_SB2_U187 ( .A(R2_SB_SB2_n752), .ZN(R2_SB_SB2_n878) );
  NOR2_X1 R2_SB_SB2_U186 ( .A1(R2_SB_SB2_n857), .A2(R2_SB_SB2_n863), .ZN(
        R2_SB_SB2_n670) );
  INV_X1 R2_SB_SB2_U185 ( .A(R2_SB_SB2_n772), .ZN(R2_SB_SB2_n883) );
  INV_X1 R2_SB_SB2_U184 ( .A(R2_SB_SB2_n618), .ZN(R2_SB_SB2_n864) );
  OAI21_X1 R2_SB_SB2_U183 ( .B1(R2_SB_SB2_n856), .B2(R2_SB_SB2_n874), .A(
        R2_SB_SB2_n893), .ZN(R2_SB_SB2_n516) );
  AOI21_X1 R2_SB_SB2_U182 ( .B1(R2_SB_SB2_n781), .B2(R2_SB_SB2_n516), .A(
        R2_SB_SB2_n515), .ZN(R2_SB_SB2_n517) );
  AOI21_X1 R2_SB_SB2_U181 ( .B1(R2_SB_SB2_n900), .B2(R2_SB_SB2_n603), .A(
        R2_SB_SB2_n783), .ZN(R2_SB_SB2_n518) );
  OAI221_X1 R2_SB_SB2_U180 ( .B1(R2_SB_SB2_n518), .B2(R2_SB_SB2_n453), .C1(
        R2_SB_SB2_n838), .C2(R2_SB_SB2_n904), .A(R2_SB_SB2_n517), .ZN(
        R2_SB_SB2_n523) );
  AOI21_X1 R2_SB_SB2_U179 ( .B1(R2_SB_SB2_n646), .B2(R2_SB_SB2_n634), .A(
        R2_SB_SB2_n633), .ZN(R2_SB_SB2_n636) );
  OAI21_X1 R2_SB_SB2_U178 ( .B1(R2_SB_SB2_n747), .B2(R2_SB_SB2_n799), .A(
        R2_SB_SB2_n882), .ZN(R2_SB_SB2_n635) );
  NAND2_X1 R2_SB_SB2_U177 ( .A1(R2_SB_SB2_n828), .A2(R2_SB_SB2_n843), .ZN(
        R2_SB_SB2_n637) );
  OAI221_X1 R2_SB_SB2_U176 ( .B1(R2_SB_SB2_n910), .B2(R2_SB_SB2_n637), .C1(
        R2_SB_SB2_n636), .C2(R2_SB_SB2_n829), .A(R2_SB_SB2_n635), .ZN(
        R2_SB_SB2_n641) );
  OAI22_X1 R2_SB_SB2_U175 ( .A1(R2_SB_SB2_n857), .A2(R2_SB_SB2_n838), .B1(
        R2_SB_SB2_n832), .B2(R2_SB_SB2_n865), .ZN(R2_SB_SB2_n469) );
  OAI21_X1 R2_SB_SB2_U174 ( .B1(R2_SB_n322), .B2(R2_SB_SB2_n845), .A(
        R2_SB_SB2_n849), .ZN(R2_SB_SB2_n471) );
  AOI221_X1 R2_SB_SB2_U173 ( .B1(R2_SB_SB2_n744), .B2(R2_SB_SB2_n471), .C1(
        R2_SB_SB2_n470), .C2(R2_SB_SB2_n863), .A(R2_SB_SB2_n469), .ZN(
        R2_SB_SB2_n476) );
  AOI221_X1 R2_SB_SB2_U172 ( .B1(R2_SB_SB2_n882), .B2(R2_SB_SB2_n792), .C1(
        R2_SB_SB2_n627), .C2(R2_SB_SB2_n702), .A(R2_SB_SB2_n698), .ZN(
        R2_SB_SB2_n583) );
  NOR2_X1 R2_SB_SB2_U171 ( .A1(R2_SB_SB2_n813), .A2(R2_SB_SB2_n694), .ZN(
        R2_SB_SB2_n695) );
  OAI221_X1 R2_SB_SB2_U170 ( .B1(R2_SB_SB2_n695), .B2(R2_SB_SB2_n851), .C1(
        R2_SB_SB2_n856), .C2(R2_SB_SB2_n878), .A(R2_SB_SB2_n904), .ZN(
        R2_SB_SB2_n697) );
  INV_X1 R2_SB_SB2_U169 ( .A(R2_SB_SB2_n801), .ZN(R2_SB_SB2_n873) );
  AOI222_X1 R2_SB_SB2_U168 ( .A1(R2_SB_SB2_n771), .A2(R2_SB_SB2_n698), .B1(
        R2_SB_SB2_n781), .B2(R2_SB_SB2_n697), .C1(R2_SB_SB2_n696), .C2(
        R2_SB_SB2_n873), .ZN(R2_SB_SB2_n741) );
  AOI22_X1 R2_SB_SB2_U167 ( .A1(R2_SB_SB2_n758), .A2(R2_SB_SB2_n694), .B1(
        R2_SB_SB2_n779), .B2(R2_SB_SB2_n863), .ZN(R2_SB_SB2_n619) );
  OAI222_X1 R2_SB_SB2_U166 ( .A1(R2_SB_SB2_n864), .A2(R2_SB_SB2_n833), .B1(
        R2_SB_n321), .B2(R2_SB_SB2_n619), .C1(R2_SB_SB2_n858), .C2(
        R2_SB_SB2_n839), .ZN(R2_SB_SB2_n620) );
  AOI221_X1 R2_SB_SB2_U165 ( .B1(R2_SB_SB2_n789), .B2(R2_SB_SB2_n628), .C1(
        R2_SB_SB2_n778), .C2(R2_SB_SB2_n771), .A(R2_SB_SB2_n620), .ZN(
        R2_SB_SB2_n621) );
  NAND2_X1 R2_SB_SB2_U164 ( .A1(R2_SB_SB2_n848), .A2(R2_SB_SB2_n841), .ZN(
        R2_SB_SB2_n616) );
  INV_X1 R2_SB_SB2_U163 ( .A(R2_SB_SB2_n615), .ZN(R2_SB_SB2_n861) );
  AOI221_X1 R2_SB_SB2_U162 ( .B1(R2_SB_SB2_n747), .B2(R2_SB_SB2_n618), .C1(
        R2_SB_SB2_n617), .C2(R2_SB_SB2_n616), .A(R2_SB_SB2_n861), .ZN(
        R2_SB_SB2_n622) );
  OAI221_X1 R2_SB_SB2_U161 ( .B1(R2_SB_SB2_n870), .B2(R2_SB_SB2_n838), .C1(
        R2_SB_SB2_n840), .C2(R2_SB_SB2_n868), .A(R2_SB_SB2_n496), .ZN(
        R2_SB_SB2_n497) );
  OAI211_X1 R2_SB_SB2_U160 ( .C1(R2_SB_SB2_n879), .C2(R2_SB_SB2_n844), .A(
        R2_SB_SB2_n711), .B(R2_SB_SB2_n491), .ZN(R2_SB_SB2_n499) );
  AOI222_X1 R2_SB_SB2_U159 ( .A1(R2_SB_SB2_n499), .A2(R2_SB_SB2_n453), .B1(
        R2_SB_SB2_n498), .B2(R2_SB_SB2_n854), .C1(R2_SB_SB2_n752), .C2(
        R2_SB_SB2_n497), .ZN(R2_SB_SB2_n527) );
  OAI222_X1 R2_SB_SB2_U158 ( .A1(R2_SB_SB2_n865), .A2(R2_SB_SB2_n838), .B1(
        R2_SB_SB2_n699), .B2(R2_SB_SB2_n868), .C1(R2_SB_n322), .C2(
        R2_SB_SB2_n858), .ZN(R2_SB_SB2_n704) );
  OAI22_X1 R2_SB_SB2_U157 ( .A1(R2_SB_SB2_n864), .A2(R2_SB_SB2_n839), .B1(
        R2_SB_SB2_n700), .B2(R2_SB_SB2_n833), .ZN(R2_SB_SB2_n701) );
  AOI222_X1 R2_SB_SB2_U156 ( .A1(R2_SB_SB2_n772), .A2(R2_SB_SB2_n704), .B1(
        R2_SB_SB2_n882), .B2(R2_SB_SB2_n703), .C1(R2_SB_SB2_n702), .C2(
        R2_SB_SB2_n701), .ZN(R2_SB_SB2_n740) );
  NOR2_X1 R2_SB_SB2_U155 ( .A1(R2_SB_SB2_n881), .A2(R2_SB_SB2_n863), .ZN(
        R2_SB_SB2_n634) );
  OAI222_X1 R2_SB_SB2_U154 ( .A1(R2_SB_n322), .A2(R2_SB_SB2_n875), .B1(
        R2_SB_SB2_n883), .B2(R2_SB_SB2_n826), .C1(R2_SB_SB2_n905), .C2(
        R2_SB_SB2_n831), .ZN(R2_SB_SB2_n707) );
  AOI211_X1 R2_SB_SB2_U153 ( .C1(R2_SB_SB2_n709), .C2(R2_SB_SB2_n708), .A(
        R2_SB_SB2_n707), .B(R2_SB_SB2_n706), .ZN(R2_SB_SB2_n710) );
  OAI222_X1 R2_SB_SB2_U152 ( .A1(R2_SB_SB2_n833), .A2(R2_SB_SB2_n898), .B1(
        R2_SB_SB2_n710), .B2(R2_SB_SB2_n859), .C1(R2_SB_SB2_n832), .C2(
        R2_SB_SB2_n800), .ZN(R2_SB_SB2_n712) );
  INV_X1 R2_SB_SB2_U151 ( .A(R2_SB_SB2_n792), .ZN(R2_SB_SB2_n845) );
  OAI221_X1 R2_SB_SB2_U150 ( .B1(R2_SB_SB2_n833), .B2(R2_SB_SB2_n774), .C1(
        R2_SB_SB2_n509), .C2(R2_SB_SB2_n829), .A(R2_SB_SB2_n508), .ZN(
        R2_SB_SB2_n510) );
  AOI221_X1 R2_SB_SB2_U149 ( .B1(R2_SB_SB2_n507), .B2(R2_SB_SB2_n506), .C1(
        R2_SB_SB2_n780), .C2(R2_SB_SB2_n684), .A(R2_SB_SB2_n505), .ZN(
        R2_SB_SB2_n512) );
  AOI221_X1 R2_SB_SB2_U148 ( .B1(R2_SB_SB2_n743), .B2(R2_SB_SB2_n684), .C1(
        R2_SB_SB2_n780), .C2(R2_SB_SB2_n627), .A(R2_SB_SB2_n510), .ZN(
        R2_SB_SB2_n511) );
  OAI222_X1 R2_SB_SB2_U147 ( .A1(R2_SB_SB2_n512), .A2(R2_SB_SB2_n905), .B1(
        R2_SB_SB2_n511), .B2(R2_SB_SB2_n883), .C1(R2_SB_SB2_n884), .C2(
        R2_SB_SB2_n844), .ZN(R2_SB_SB2_n513) );
  INV_X1 R2_SB_SB2_U146 ( .A(R2_SB_SB2_n659), .ZN(R2_SB_SB2_n867) );
  AOI221_X1 R2_SB_SB2_U145 ( .B1(R2_SB_SB2_n794), .B2(R2_SB_SB2_n730), .C1(
        R2_SB_SB2_n742), .C2(R2_SB_SB2_n780), .A(R2_SB_SB2_n867), .ZN(
        R2_SB_SB2_n574) );
  NOR4_X1 R2_SB_SB2_U144 ( .A1(R2_SB_SB2_n452), .A2(R2_SB_SB2_n872), .A3(
        R2_SB_SB2_n849), .A4(R2_SB_SB2_n862), .ZN(R2_SB_SB2_n640) );
  NOR2_X1 R2_SB_SB2_U143 ( .A1(R2_SB_SB2_n89), .A2(R2_SB_SB2_n843), .ZN(
        R2_SB_SB2_n603) );
  NOR2_X1 R2_SB_SB2_U142 ( .A1(R2_SB_SB2_n872), .A2(R2_SB_SB2_n863), .ZN(
        R2_SB_SB2_n812) );
  NOR2_X1 R2_SB_SB2_U141 ( .A1(R2_SB_SB2_n863), .A2(R2_SB_SB2_n854), .ZN(
        R2_SB_SB2_n507) );
  AOI222_X1 R2_SB_SB2_U140 ( .A1(R2_SB_SB2_n782), .A2(R2_SB_SB2_n781), .B1(
        R2_SB_SB2_n780), .B2(R2_SB_SB2_n779), .C1(R2_SB_SB2_n778), .C2(
        R2_SB_SB2_n791), .ZN(R2_SB_SB2_n784) );
  INV_X1 R2_SB_SB2_U139 ( .A(R2_SB_SB2_n795), .ZN(R2_SB_SB2_n838) );
  AOI22_X1 R2_SB_SB2_U138 ( .A1(R2_SB_SB2_n724), .A2(R2_SB_SB2_n810), .B1(
        R2_SB_SB2_n744), .B2(R2_SB_SB2_n723), .ZN(R2_SB_SB2_n726) );
  INV_X1 R2_SB_SB2_U137 ( .A(R2_SB_SB2_n722), .ZN(R2_SB_SB2_n896) );
  INV_X1 R2_SB_SB2_U136 ( .A(R2_SB_SB2_n725), .ZN(R2_SB_SB2_n846) );
  OAI222_X1 R2_SB_SB2_U135 ( .A1(R2_SB_SB2_n849), .A2(R2_SB_SB2_n896), .B1(
        R2_SB_SB2_n726), .B2(R2_SB_SB2_n878), .C1(R2_SB_SB2_n846), .C2(
        R2_SB_SB2_n910), .ZN(R2_SB_SB2_n735) );
  OAI222_X1 R2_SB_SB2_U134 ( .A1(R2_SB_SB2_n853), .A2(R2_SB_SB2_n829), .B1(
        R2_SB_SB2_n608), .B2(R2_SB_SB2_n826), .C1(R2_SB_SB2_n870), .C2(
        R2_SB_SB2_n831), .ZN(R2_SB_SB2_n465) );
  NOR3_X1 R2_SB_SB2_U133 ( .A1(R2_SB_SB2_n877), .A2(R2_SB_SB2_n638), .A3(
        R2_SB_SB2_n679), .ZN(R2_SB_SB2_n466) );
  INV_X1 R2_SB_SB2_U132 ( .A(R2_SB_SB2_n465), .ZN(R2_SB_SB2_n871) );
  OAI222_X1 R2_SB_SB2_U131 ( .A1(R2_SB_SB2_n871), .A2(R2_SB_SB2_n883), .B1(
        R2_SB_SB2_n849), .B2(R2_SB_SB2_n769), .C1(R2_SB_SB2_n466), .C2(
        R2_SB_SB2_n834), .ZN(R2_SB_SB2_n484) );
  INV_X1 R2_SB_SB2_U130 ( .A(R2_SB_SB2_n782), .ZN(R2_SB_SB2_n849) );
  NOR2_X1 R2_SB_SB2_U129 ( .A1(R2_SB_SB2_n830), .A2(R2_SB_SB2_n854), .ZN(
        R2_SB_SB2_n627) );
  NOR2_X1 R2_SB_SB2_U128 ( .A1(R2_SB_SB2_n881), .A2(R2_SB_SB2_n872), .ZN(
        R2_SB_SB2_n669) );
  INV_X1 R2_SB_SB2_U127 ( .A(R2_SB_SB2_n702), .ZN(R2_SB_SB2_n905) );
  NOR2_X1 R2_SB_SB2_U126 ( .A1(R2_SB_SB2_n453), .A2(R2_SB_SB2_n830), .ZN(
        R2_SB_SB2_n766) );
  NOR3_X1 R2_SB_SB2_U125 ( .A1(R2_SB_SB2_n828), .A2(R2_SB_SB2_n854), .A3(
        R2_SB_SB2_n908), .ZN(R2_SB_SB2_n673) );
  NOR2_X1 R2_SB_SB2_U124 ( .A1(R2_SB_SB2_n89), .A2(R2_SB_SB2_n830), .ZN(
        R2_SB_SB2_n771) );
  NOR2_X1 R2_SB_SB2_U123 ( .A1(R2_SB_SB2_n863), .A2(R2_SB_SB2_n843), .ZN(
        R2_SB_SB2_n778) );
  NOR2_X1 R2_SB_SB2_U122 ( .A1(R2_SB_SB2_n830), .A2(R2_SB_n322), .ZN(
        R2_SB_SB2_n779) );
  AOI21_X1 R2_SB_SB2_U121 ( .B1(R2_SB_SB2_n826), .B2(R2_SB_SB2_n833), .A(
        R2_SB_SB2_n800), .ZN(R2_SB_SB2_n549) );
  INV_X1 R2_SB_SB2_U120 ( .A(R2_SB_SB2_n549), .ZN(R2_SB_SB2_n902) );
  AND3_X1 R2_SB_SB2_U119 ( .A1(R2_SB_SB2_n548), .A2(R2_SB_SB2_n838), .A3(
        R2_SB_SB2_n849), .ZN(R2_SB_SB2_n550) );
  OR3_X1 R2_SB_SB2_U118 ( .A1(R2_SB_SB2_n864), .A2(R2_SB_SB2_n814), .A3(
        R2_SB_SB2_n890), .ZN(R2_SB_SB2_n815) );
  INV_X1 R2_SB_SB2_U117 ( .A(R2_SB_SB2_n519), .ZN(R2_SB_SB2_n886) );
  INV_X1 R2_SB_SB2_U116 ( .A(R2_SB_SB2_n790), .ZN(R2_SB_SB2_n866) );
  NAND2_X1 R2_SB_SB2_U115 ( .A1(R2_SB_SB2_n874), .A2(R2_SB_SB2_n901), .ZN(
        R2_SB_SB2_n728) );
  NAND2_X1 R2_SB_SB2_U114 ( .A1(R2_SB_SB2_n890), .A2(R2_SB_SB2_n874), .ZN(
        R2_SB_SB2_n536) );
  NAND2_X1 R2_SB_SB2_U113 ( .A1(R2_SB_SB2_n836), .A2(R2_SB_SB2_n826), .ZN(
        R2_SB_SB2_n723) );
  NAND2_X1 R2_SB_SB2_U112 ( .A1(R2_SB_SB2_n905), .A2(R2_SB_SB2_n875), .ZN(
        R2_SB_SB2_n589) );
  INV_X1 R2_SB_SB2_U111 ( .A(R2_SB_SB2_n627), .ZN(R2_SB_SB2_n856) );
  NAND2_X1 R2_SB_SB2_U110 ( .A1(R2_SB_SB2_n836), .A2(R2_SB_SB2_n829), .ZN(
        R2_SB_SB2_n748) );
  AND2_X1 R2_SB_SB2_U109 ( .A1(R2_SB_SB2_n766), .A2(R2_SB_SB2_n671), .ZN(
        R2_SB_SB2_n555) );
  INV_X1 R2_SB_SB2_U108 ( .A(R2_SB_SB2_n812), .ZN(R2_SB_SB2_n875) );
  OAI21_X1 R2_SB_SB2_U107 ( .B1(R2_SB_SB2_n847), .B2(R2_SB_SB2_n895), .A(
        R2_SB_SB2_n800), .ZN(R2_SB_SB2_n806) );
  NAND2_X1 R2_SB_SB2_U106 ( .A1(R2_SB_SB2_n628), .A2(R2_SB_SB2_n634), .ZN(
        R2_SB_SB2_n769) );
  NAND2_X1 R2_SB_SB2_U105 ( .A1(R2_SB_SB2_n507), .A2(R2_SB_SB2_n669), .ZN(
        R2_SB_SB2_n588) );
  INV_X1 R2_SB_SB2_U104 ( .A(R2_SB_SB2_n634), .ZN(R2_SB_SB2_n903) );
  INV_X1 R2_SB_SB2_U103 ( .A(R2_SB_SB2_n778), .ZN(R2_SB_SB2_n865) );
  NOR2_X1 R2_SB_SB2_U102 ( .A1(R2_SB_SB2_n730), .A2(R2_SB_SB2_n758), .ZN(
        R2_SB_SB2_n685) );
  AOI21_X1 R2_SB_SB2_U101 ( .B1(R2_SB_SB2_n588), .B2(R2_SB_SB2_n773), .A(
        R2_SB_SB2_n836), .ZN(R2_SB_SB2_n460) );
  AOI21_X1 R2_SB_SB2_U100 ( .B1(R2_SB_SB2_n802), .B2(R2_SB_SB2_n801), .A(
        R2_SB_SB2_n835), .ZN(R2_SB_SB2_n803) );
  INV_X1 R2_SB_SB2_U99 ( .A(R2_SB_SB2_n672), .ZN(R2_SB_SB2_n888) );
  NOR4_X1 R2_SB_SB2_U98 ( .A1(R2_SB_SB2_n675), .A2(R2_SB_SB2_n888), .A3(
        R2_SB_SB2_n674), .A4(R2_SB_SB2_n673), .ZN(R2_SB_SB2_n676) );
  NAND2_X1 R2_SB_SB2_U97 ( .A1(R2_SB_SB2_n778), .A2(R2_SB_SB2_n669), .ZN(
        R2_SB_SB2_n573) );
  INV_X1 R2_SB_SB2_U96 ( .A(R2_SB_SB2_n648), .ZN(R2_SB_SB2_n882) );
  NOR2_X1 R2_SB_SB2_U95 ( .A1(R2_SB_SB2_n849), .A2(R2_SB_SB2_n89), .ZN(
        R2_SB_SB2_n502) );
  NOR2_X1 R2_SB_SB2_U94 ( .A1(R2_SB_SB2_n851), .A2(R2_SB_n322), .ZN(
        R2_SB_SB2_n470) );
  NOR2_X1 R2_SB_SB2_U93 ( .A1(R2_SB_SB2_n853), .A2(R2_SB_SB2_n903), .ZN(
        R2_SB_SB2_n514) );
  INV_X1 R2_SB_SB2_U92 ( .A(R2_SB_SB2_n604), .ZN(R2_SB_SB2_n844) );
  NOR2_X1 R2_SB_SB2_U91 ( .A1(R2_SB_SB2_n862), .A2(R2_SB_SB2_n883), .ZN(
        R2_SB_SB2_n534) );
  INV_X1 R2_SB_SB2_U90 ( .A(R2_SB_SB2_n603), .ZN(R2_SB_SB2_n848) );
  INV_X1 R2_SB_SB2_U89 ( .A(R2_SB_SB2_n802), .ZN(R2_SB_SB2_n877) );
  NOR2_X1 R2_SB_SB2_U88 ( .A1(R2_SB_SB2_n905), .A2(R2_SB_SB2_n866), .ZN(
        R2_SB_SB2_n671) );
  OAI22_X1 R2_SB_SB2_U87 ( .A1(R2_SB_SB2_n730), .A2(R2_SB_SB2_n905), .B1(
        R2_SB_SB2_n901), .B2(R2_SB_SB2_n851), .ZN(R2_SB_SB2_n462) );
  OAI22_X1 R2_SB_SB2_U86 ( .A1(R2_SB_SB2_n875), .A2(R2_SB_SB2_n833), .B1(
        R2_SB_SB2_n874), .B2(R2_SB_SB2_n832), .ZN(R2_SB_SB2_n804) );
  OAI22_X1 R2_SB_SB2_U85 ( .A1(R2_SB_SB2_n665), .A2(R2_SB_SB2_n892), .B1(
        R2_SB_SB2_n841), .B2(R2_SB_SB2_n801), .ZN(R2_SB_SB2_n666) );
  INV_X1 R2_SB_SB2_U84 ( .A(R2_SB_SB2_n758), .ZN(R2_SB_SB2_n847) );
  AOI21_X1 R2_SB_SB2_U83 ( .B1(R2_SB_SB2_n868), .B2(R2_SB_SB2_n845), .A(
        R2_SB_SB2_n785), .ZN(R2_SB_SB2_n687) );
  OAI22_X1 R2_SB_SB2_U82 ( .A1(R2_SB_SB2_n831), .A2(R2_SB_SB2_n895), .B1(
        R2_SB_n321), .B2(R2_SB_SB2_n648), .ZN(R2_SB_SB2_n532) );
  AOI22_X1 R2_SB_SB2_U81 ( .A1(R2_SB_SB2_n758), .A2(R2_SB_n322), .B1(
        R2_SB_SB2_n771), .B2(R2_SB_SB2_n452), .ZN(R2_SB_SB2_n699) );
  INV_X1 R2_SB_SB2_U80 ( .A(R2_SB_SB2_n771), .ZN(R2_SB_SB2_n831) );
  NOR2_X1 R2_SB_SB2_U79 ( .A1(R2_SB_SB2_n842), .A2(R2_SB_SB2_n898), .ZN(
        R2_SB_SB2_n675) );
  NOR2_X1 R2_SB_SB2_U78 ( .A1(R2_SB_SB2_n868), .A2(R2_SB_SB2_n890), .ZN(
        R2_SB_SB2_n576) );
  NOR2_X1 R2_SB_SB2_U77 ( .A1(R2_SB_SB2_n774), .A2(R2_SB_SB2_n890), .ZN(
        R2_SB_SB2_n565) );
  NOR2_X1 R2_SB_SB2_U76 ( .A1(R2_SB_SB2_n845), .A2(R2_SB_SB2_n89), .ZN(
        R2_SB_SB2_n725) );
  NOR2_X1 R2_SB_SB2_U75 ( .A1(R2_SB_SB2_n853), .A2(R2_SB_SB2_n890), .ZN(
        R2_SB_SB2_n633) );
  NOR2_X1 R2_SB_SB2_U74 ( .A1(R2_SB_SB2_n868), .A2(R2_SB_SB2_n905), .ZN(
        R2_SB_SB2_n754) );
  NOR2_X1 R2_SB_SB2_U73 ( .A1(R2_SB_SB2_n869), .A2(R2_SB_SB2_n905), .ZN(
        R2_SB_SB2_n698) );
  NOR2_X1 R2_SB_SB2_U72 ( .A1(R2_SB_SB2_n898), .A2(R2_SB_SB2_n845), .ZN(
        R2_SB_SB2_n756) );
  NOR2_X1 R2_SB_SB2_U71 ( .A1(R2_SB_SB2_n774), .A2(R2_SB_SB2_n905), .ZN(
        R2_SB_SB2_n638) );
  NOR2_X1 R2_SB_SB2_U70 ( .A1(R2_SB_SB2_n870), .A2(R2_SB_SB2_n890), .ZN(
        R2_SB_SB2_n727) );
  OAI22_X1 R2_SB_SB2_U69 ( .A1(R2_SB_SB2_n453), .A2(R2_SB_SB2_n879), .B1(
        R2_SB_SB2_n89), .B2(R2_SB_SB2_n880), .ZN(R2_SB_SB2_n538) );
  AOI211_X1 R2_SB_SB2_U68 ( .C1(R2_SB_SB2_n576), .C2(R2_SB_SB2_n89), .A(
        R2_SB_SB2_n538), .B(R2_SB_SB2_n722), .ZN(R2_SB_SB2_n543) );
  INV_X1 R2_SB_SB2_U67 ( .A(R2_SB_SB2_n779), .ZN(R2_SB_SB2_n833) );
  NOR3_X1 R2_SB_SB2_U66 ( .A1(R2_SB_SB2_n841), .A2(R2_SB_SB2_n858), .A3(
        R2_SB_SB2_n874), .ZN(R2_SB_SB2_n521) );
  INV_X1 R2_SB_SB2_U65 ( .A(R2_SB_SB2_n766), .ZN(R2_SB_SB2_n835) );
  NOR2_X1 R2_SB_SB2_U64 ( .A1(R2_SB_SB2_n838), .A2(R2_SB_SB2_n453), .ZN(
        R2_SB_SB2_n742) );
  INV_X1 R2_SB_SB2_U63 ( .A(R2_SB_SB2_n730), .ZN(R2_SB_SB2_n858) );
  NOR2_X1 R2_SB_SB2_U62 ( .A1(R2_SB_SB2_n878), .A2(R2_SB_SB2_n869), .ZN(
        R2_SB_SB2_n713) );
  NOR2_X1 R2_SB_SB2_U61 ( .A1(R2_SB_SB2_n833), .A2(R2_SB_SB2_n453), .ZN(
        R2_SB_SB2_n799) );
  AOI22_X1 R2_SB_SB2_U60 ( .A1(R2_SB_SB2_n877), .A2(R2_SB_SB2_n452), .B1(
        R2_SB_SB2_n781), .B2(R2_SB_SB2_n669), .ZN(R2_SB_SB2_n500) );
  OAI211_X1 R2_SB_SB2_U59 ( .C1(R2_SB_SB2_n89), .C2(R2_SB_SB2_n893), .A(
        R2_SB_SB2_n907), .B(R2_SB_SB2_n500), .ZN(R2_SB_SB2_n501) );
  AOI222_X1 R2_SB_SB2_U58 ( .A1(R2_SB_SB2_n591), .A2(R2_SB_SB2_n748), .B1(
        R2_SB_SB2_n502), .B2(R2_SB_SB2_n679), .C1(R2_SB_SB2_n758), .C2(
        R2_SB_SB2_n501), .ZN(R2_SB_SB2_n526) );
  OAI222_X1 R2_SB_SB2_U57 ( .A1(R2_SB_SB2_n845), .A2(R2_SB_SB2_n880), .B1(
        R2_SB_SB2_n835), .B2(R2_SB_SB2_n898), .C1(R2_SB_SB2_n836), .C2(
        R2_SB_SB2_n894), .ZN(R2_SB_SB2_n602) );
  NOR2_X1 R2_SB_SB2_U56 ( .A1(R2_SB_SB2_n883), .A2(R2_SB_SB2_n869), .ZN(
        R2_SB_SB2_n755) );
  NOR2_X1 R2_SB_SB2_U55 ( .A1(R2_SB_SB2_n862), .A2(R2_SB_SB2_n890), .ZN(
        R2_SB_SB2_n753) );
  NOR2_X1 R2_SB_SB2_U54 ( .A1(R2_SB_SB2_n862), .A2(R2_SB_SB2_n905), .ZN(
        R2_SB_SB2_n759) );
  NOR2_X1 R2_SB_SB2_U53 ( .A1(R2_SB_SB2_n862), .A2(R2_SB_SB2_n878), .ZN(
        R2_SB_SB2_n591) );
  NOR2_X1 R2_SB_SB2_U52 ( .A1(R2_SB_SB2_n869), .A2(R2_SB_SB2_n890), .ZN(
        R2_SB_SB2_n679) );
  INV_X1 R2_SB_SB2_U51 ( .A(R2_SB_SB2_n669), .ZN(R2_SB_SB2_n890) );
  NOR2_X2 R2_SB_SB2_U50 ( .A1(R2_SB_SB2_n89), .A2(R2_SB_SB2_n453), .ZN(
        R2_SB_SB2_n781) );
  NOR2_X2 R2_SB_SB2_U49 ( .A1(R2_SB_SB2_n89), .A2(R2_SB_SB2_n452), .ZN(
        R2_SB_SB2_n684) );
  NOR3_X1 R2_SB_SB2_U48 ( .A1(R2_SB_SB2_n878), .A2(R2_SB_SB2_n866), .A3(
        R2_SB_SB2_n838), .ZN(R2_SB_SB2_n674) );
  NOR2_X1 R2_SB_SB2_U47 ( .A1(R2_SB_SB2_n840), .A2(R2_SB_SB2_n452), .ZN(
        R2_SB_SB2_n747) );
  NOR2_X1 R2_SB_SB2_U46 ( .A1(R2_SB_SB2_n453), .A2(R2_SB_n322), .ZN(
        R2_SB_SB2_n810) );
  INV_X1 R2_SB_SB2_U45 ( .A(R2_SB_SB2_n633), .ZN(R2_SB_SB2_n891) );
  INV_X1 R2_SB_SB2_U44 ( .A(R2_SB_SB2_n534), .ZN(R2_SB_SB2_n885) );
  INV_X1 R2_SB_SB2_U43 ( .A(R2_SB_SB2_n470), .ZN(R2_SB_SB2_n852) );
  INV_X1 R2_SB_SB2_U42 ( .A(R2_SB_SB2_n502), .ZN(R2_SB_SB2_n850) );
  INV_X1 R2_SB_SB2_U41 ( .A(R2_SB_SB2_n514), .ZN(R2_SB_SB2_n904) );
  INV_X1 R2_SB_SB2_U40 ( .A(R2_SB_SB2_n698), .ZN(R2_SB_SB2_n906) );
  INV_X1 R2_SB_SB2_U39 ( .A(R2_SB_SB2_n638), .ZN(R2_SB_SB2_n908) );
  INV_X1 R2_SB_SB2_U38 ( .A(R2_SB_SB2_n565), .ZN(R2_SB_SB2_n892) );
  INV_X1 R2_SB_SB2_U37 ( .A(R2_SB_SB2_n753), .ZN(R2_SB_SB2_n893) );
  INV_X1 R2_SB_SB2_U36 ( .A(R2_SB_SB2_n727), .ZN(R2_SB_SB2_n894) );
  INV_X1 R2_SB_SB2_U35 ( .A(R2_SB_SB2_n755), .ZN(R2_SB_SB2_n884) );
  INV_X1 R2_SB_SB2_U34 ( .A(R2_SB_SB2_n799), .ZN(R2_SB_SB2_n834) );
  NAND2_X1 R2_SB_SB2_U33 ( .A1(R2_SB_SB2_n781), .A2(R2_SB_SB2_n671), .ZN(
        R2_SB_SB2_n716) );
  INV_X1 R2_SB_SB2_U32 ( .A(R2_SB_SB2_n588), .ZN(R2_SB_SB2_n900) );
  INV_X1 R2_SB_SB2_U31 ( .A(R2_SB_SB2_n759), .ZN(R2_SB_SB2_n907) );
  INV_X1 R2_SB_SB2_U30 ( .A(R2_SB_SB2_n747), .ZN(R2_SB_SB2_n841) );
  INV_X1 R2_SB_SB2_U29 ( .A(R2_SB_SB2_n713), .ZN(R2_SB_SB2_n879) );
  INV_X1 R2_SB_SB2_U28 ( .A(R2_SB_SB2_n591), .ZN(R2_SB_SB2_n880) );
  INV_X1 R2_SB_SB2_U27 ( .A(R2_SB_SB2_n742), .ZN(R2_SB_SB2_n839) );
  AOI21_X1 R2_SB_SB2_U26 ( .B1(R2_SB_SB2_n848), .B2(R2_SB_SB2_n852), .A(
        R2_SB_SB2_n910), .ZN(R2_SB_SB2_n461) );
  AOI21_X1 R2_SB_SB2_U25 ( .B1(R2_SB_SB2_n831), .B2(R2_SB_SB2_n835), .A(
        R2_SB_SB2_n890), .ZN(R2_SB_SB2_n796) );
  INV_X1 R2_SB_SB2_U24 ( .A(R2_SB_SB2_n684), .ZN(R2_SB_SB2_n827) );
  AOI22_X1 R2_SB_SB2_U23 ( .A1(R2_SB_SB2_n877), .A2(R2_SB_n322), .B1(
        R2_SB_SB2_n713), .B2(R2_SB_SB2_n828), .ZN(R2_SB_SB2_n649) );
  INV_X1 R2_SB_SB2_U22 ( .A(R2_SB_SB2_n754), .ZN(R2_SB_SB2_n910) );
  INV_X1 R2_SB_SB2_U21 ( .A(R2_SB_SB2_n781), .ZN(R2_SB_SB2_n828) );
  INV_X1 R2_SB_SB2_U20 ( .A(R2_SB_SB2_n576), .ZN(R2_SB_SB2_n898) );
  INV_X1 R2_SB_SB2_U19 ( .A(R2_SB_SB2_n679), .ZN(R2_SB_SB2_n895) );
  NOR2_X1 R2_SB_SB2_U18 ( .A1(R2_SB_SB2_n831), .A2(R2_SB_SB2_n452), .ZN(
        R2_SB_SB2_n708) );
  OAI221_X1 R2_SB_SB2_U17 ( .B1(R2_SB_n322), .B2(R2_SB_SB2_n906), .C1(
        R2_SB_SB2_n890), .C2(R2_SB_SB2_n826), .A(R2_SB_SB2_n769), .ZN(
        R2_SB_SB2_n590) );
  NOR2_X1 R2_SB_SB2_U16 ( .A1(R2_SB_SB2_n895), .A2(R2_SB_SB2_n452), .ZN(
        R2_SB_SB2_n722) );
  INV_X1 R2_SB_SB2_U15 ( .A(R2_SB_SB2_n810), .ZN(R2_SB_SB2_n829) );
  NOR2_X1 R2_SB_SB2_U14 ( .A1(R2_SB_n321), .A2(R2_SB_n322), .ZN(R2_SB_SB2_n628) );
  INV_X1 R2_SB_SB2_U13 ( .A(R2_SB_SB2_n708), .ZN(R2_SB_SB2_n832) );
  INV_X1 R2_SB_SB2_U12 ( .A(R2_SB_SB2_n628), .ZN(R2_SB_SB2_n826) );
  NOR2_X1 R2_SB_SB2_U11 ( .A1(R2_SB_SB2_n863), .A2(R2_SB_n325), .ZN(
        R2_SB_SB2_n744) );
  NOR2_X1 R2_SB_SB2_U10 ( .A1(R2_SB_SB2_n881), .A2(R2_SB_n327), .ZN(
        R2_SB_SB2_n772) );
  NOR2_X1 R2_SB_SB2_U9 ( .A1(R2_SB_SB2_n89), .A2(R2_SB_n323), .ZN(
        R2_SB_SB2_n791) );
  NOR2_X1 R2_SB_SB2_U8 ( .A1(R2_SB_SB2_n872), .A2(R2_SB_n328), .ZN(
        R2_SB_SB2_n752) );
  NOR2_X1 R2_SB_SB2_U7 ( .A1(R2_SB_SB2_n854), .A2(R2_SB_SB2_n843), .ZN(
        R2_SB_SB2_n730) );
  NOR2_X1 R2_SB_SB2_U6 ( .A1(R2_SB_SB2_n843), .A2(R2_SB_n326), .ZN(
        R2_SB_SB2_n780) );
  NOR2_X1 R2_SB_SB2_U5 ( .A1(R2_SB_n323), .A2(R2_SB_n324), .ZN(R2_SB_SB2_n743)
         );
  INV_X1 R2_SB_SB2_U4 ( .A(R2_SB_n324), .ZN(R2_SB_SB2_n843) );
  NOR2_X1 R2_SB_SB2_U3 ( .A1(R2_SB_SB2_n453), .A2(R2_SB_n323), .ZN(
        R2_SB_SB2_n696) );
  NOR2_X1 R2_SB_SB2_U2 ( .A1(R2_SB_SB2_n881), .A2(R2_SB_n326), .ZN(
        R2_SB_SB2_n798) );
  NOR2_X1 R2_SB_SB2_U1 ( .A1(R2_SB_SB2_n843), .A2(R2_SB_n325), .ZN(
        R2_SB_SB2_n789) );
  NAND3_X1 R2_SB_SB2_U464 ( .A1(R2_SB_SB2_n772), .A2(R2_SB_SB2_n670), .A3(
        R2_SB_SB2_n794), .ZN(R2_SB_SB2_n519) );
  OAI33_X1 R2_SB_SB2_U463 ( .A1(R2_SB_SB2_n838), .A2(R2_SB_SB2_n858), .A3(
        R2_SB_SB2_n905), .B1(R2_SB_SB2_n853), .B2(R2_SB_SB2_n830), .B3(
        R2_SB_SB2_n874), .ZN(R2_SB_SB2_n467) );
  NAND3_X1 R2_SB_SB2_U462 ( .A1(R2_SB_SB2_n507), .A2(R2_SB_SB2_n702), .A3(
        R2_SB_SB2_n758), .ZN(R2_SB_SB2_n677) );
  OAI33_X1 R2_SB_SB2_U461 ( .A1(R2_SB_SB2_n828), .A2(R2_SB_n328), .A3(
        R2_SB_n323), .B1(R2_SB_SB2_n472), .B2(R2_SB_SB2_n854), .B3(
        R2_SB_SB2_n829), .ZN(R2_SB_SB2_n473) );
  NAND4_X1 R2_SB_SB2_U460 ( .A1(R2_SB_SB2_n488), .A2(R2_SB_SB2_n487), .A3(
        R2_SB_SB2_n486), .A4(R2_SB_SB2_n485), .ZN(R2_SB_n313) );
  NAND3_X1 R2_SB_SB2_U459 ( .A1(R2_SB_SB2_n781), .A2(R2_SB_n323), .A3(
        R2_SB_SB2_n798), .ZN(R2_SB_SB2_n494) );
  NAND4_X1 R2_SB_SB2_U458 ( .A1(R2_SB_SB2_n743), .A2(R2_SB_SB2_n628), .A3(
        R2_SB_SB2_n767), .A4(R2_SB_n328), .ZN(R2_SB_SB2_n493) );
  NAND3_X1 R2_SB_SB2_U457 ( .A1(R2_SB_SB2_n813), .A2(R2_SB_SB2_n830), .A3(
        R2_SB_SB2_n684), .ZN(R2_SB_SB2_n492) );
  NAND3_X1 R2_SB_SB2_U456 ( .A1(R2_SB_SB2_n494), .A2(R2_SB_SB2_n493), .A3(
        R2_SB_SB2_n492), .ZN(R2_SB_SB2_n498) );
  NAND3_X1 R2_SB_SB2_U455 ( .A1(R2_SB_SB2_n844), .A2(R2_SB_SB2_n836), .A3(
        R2_SB_SB2_n548), .ZN(R2_SB_SB2_n506) );
  OAI33_X1 R2_SB_SB2_U454 ( .A1(R2_SB_SB2_n827), .A2(R2_SB_SB2_n856), .A3(
        R2_SB_SB2_n903), .B1(R2_SB_SB2_n898), .B2(R2_SB_SB2_n843), .B3(
        R2_SB_SB2_n826), .ZN(R2_SB_SB2_n515) );
  NAND3_X1 R2_SB_SB2_U453 ( .A1(R2_SB_SB2_n671), .A2(R2_SB_SB2_n453), .A3(
        R2_SB_n323), .ZN(R2_SB_SB2_n816) );
  NAND3_X1 R2_SB_SB2_U452 ( .A1(R2_SB_SB2_n670), .A2(R2_SB_SB2_n669), .A3(
        R2_SB_SB2_n779), .ZN(R2_SB_SB2_n672) );
  NAND3_X1 R2_SB_SB2_U451 ( .A1(R2_SB_SB2_n816), .A2(R2_SB_SB2_n519), .A3(
        R2_SB_SB2_n672), .ZN(R2_SB_SB2_n522) );
  OAI33_X1 R2_SB_SB2_U450 ( .A1(R2_SB_SB2_n832), .A2(R2_SB_SB2_n864), .A3(
        R2_SB_SB2_n890), .B1(R2_SB_SB2_n829), .B2(R2_SB_n328), .B3(
        R2_SB_SB2_n866), .ZN(R2_SB_SB2_n520) );
  NAND4_X1 R2_SB_SB2_U449 ( .A1(R2_SB_SB2_n527), .A2(R2_SB_SB2_n526), .A3(
        R2_SB_SB2_n525), .A4(R2_SB_SB2_n524), .ZN(R2_SB_n314) );
  NAND3_X1 R2_SB_SB2_U448 ( .A1(R2_SB_SB2_n744), .A2(R2_SB_SB2_n603), .A3(
        R2_SB_SB2_n696), .ZN(R2_SB_SB2_n546) );
  NAND3_X1 R2_SB_SB2_U447 ( .A1(R2_SB_SB2_n684), .A2(R2_SB_SB2_n854), .A3(
        R2_SB_SB2_n709), .ZN(R2_SB_SB2_n582) );
  OAI33_X1 R2_SB_SB2_U446 ( .A1(R2_SB_SB2_n859), .A2(R2_SB_SB2_n830), .A3(
        R2_SB_SB2_n901), .B1(R2_SB_SB2_n876), .B2(R2_SB_n322), .B3(
        R2_SB_SB2_n685), .ZN(R2_SB_SB2_n557) );
  NAND4_X1 R2_SB_SB2_U445 ( .A1(R2_SB_SB2_n561), .A2(R2_SB_SB2_n560), .A3(
        R2_SB_SB2_n559), .A4(R2_SB_SB2_n558), .ZN(R2_SB_n315) );
  NAND3_X1 R2_SB_SB2_U444 ( .A1(R2_SB_SB2_n830), .A2(R2_SB_SB2_n872), .A3(
        R2_SB_SB2_n709), .ZN(R2_SB_SB2_n566) );
  NAND4_X1 R2_SB_SB2_U443 ( .A1(R2_SB_SB2_n566), .A2(R2_SB_SB2_n894), .A3(
        R2_SB_SB2_n800), .A4(R2_SB_SB2_n648), .ZN(R2_SB_SB2_n569) );
  NAND3_X1 R2_SB_SB2_U442 ( .A1(R2_SB_n321), .A2(R2_SB_n324), .A3(
        R2_SB_SB2_n744), .ZN(R2_SB_SB2_n659) );
  NAND3_X1 R2_SB_SB2_U441 ( .A1(R2_SB_SB2_n758), .A2(R2_SB_SB2_n854), .A3(
        R2_SB_SB2_n709), .ZN(R2_SB_SB2_n587) );
  NAND3_X1 R2_SB_SB2_U440 ( .A1(R2_SB_SB2_n743), .A2(R2_SB_n321), .A3(
        R2_SB_SB2_n882), .ZN(R2_SB_SB2_n592) );
  NAND4_X1 R2_SB_SB2_U439 ( .A1(R2_SB_SB2_n601), .A2(R2_SB_SB2_n600), .A3(
        R2_SB_SB2_n599), .A4(R2_SB_SB2_n598), .ZN(R2_SB_n316) );
  NAND4_X1 R2_SB_SB2_U438 ( .A1(R2_SB_SB2_n645), .A2(R2_SB_SB2_n644), .A3(
        R2_SB_SB2_n643), .A4(R2_SB_SB2_n642), .ZN(R2_SB_n317) );
  NAND3_X1 R2_SB_SB2_U437 ( .A1(R2_SB_SB2_n684), .A2(R2_SB_SB2_n843), .A3(
        R2_SB_SB2_n744), .ZN(R2_SB_SB2_n660) );
  NAND3_X1 R2_SB_SB2_U436 ( .A1(R2_SB_n321), .A2(R2_SB_SB2_n854), .A3(
        R2_SB_SB2_n792), .ZN(R2_SB_SB2_n658) );
  NAND4_X1 R2_SB_SB2_U435 ( .A1(R2_SB_SB2_n660), .A2(R2_SB_SB2_n659), .A3(
        R2_SB_SB2_n658), .A4(R2_SB_SB2_n657), .ZN(R2_SB_SB2_n668) );
  OAI33_X1 R2_SB_SB2_U434 ( .A1(R2_SB_SB2_n862), .A2(R2_SB_n328), .A3(
        R2_SB_SB2_n847), .B1(R2_SB_SB2_n903), .B2(R2_SB_SB2_n858), .B3(
        R2_SB_SB2_n830), .ZN(R2_SB_SB2_n661) );
  NAND3_X1 R2_SB_SB2_U433 ( .A1(R2_SB_SB2_n670), .A2(R2_SB_SB2_n669), .A3(
        R2_SB_SB2_n766), .ZN(R2_SB_SB2_n717) );
  NAND4_X1 R2_SB_SB2_U432 ( .A1(R2_SB_SB2_n717), .A2(R2_SB_SB2_n716), .A3(
        R2_SB_SB2_n677), .A4(R2_SB_SB2_n676), .ZN(R2_SB_SB2_n689) );
  OAI33_X1 R2_SB_SB2_U431 ( .A1(R2_SB_SB2_n839), .A2(R2_SB_SB2_n870), .A3(
        R2_SB_SB2_n883), .B1(R2_SB_SB2_n827), .B2(R2_SB_SB2_n685), .B3(
        R2_SB_SB2_n903), .ZN(R2_SB_SB2_n686) );
  NAND4_X1 R2_SB_SB2_U430 ( .A1(R2_SB_SB2_n693), .A2(R2_SB_SB2_n692), .A3(
        R2_SB_SB2_n691), .A4(R2_SB_SB2_n690), .ZN(R2_SB_n318) );
  NAND3_X1 R2_SB_SB2_U429 ( .A1(R2_SB_SB2_n845), .A2(R2_SB_SB2_n838), .A3(
        R2_SB_SB2_n829), .ZN(R2_SB_SB2_n703) );
  OAI33_X1 R2_SB_SB2_U428 ( .A1(R2_SB_SB2_n876), .A2(R2_SB_n321), .A3(
        R2_SB_SB2_n830), .B1(R2_SB_SB2_n705), .B2(R2_SB_SB2_n835), .B3(
        R2_SB_SB2_n901), .ZN(R2_SB_SB2_n706) );
  NAND3_X1 R2_SB_SB2_U427 ( .A1(R2_SB_n325), .A2(R2_SB_SB2_n714), .A3(
        R2_SB_n328), .ZN(R2_SB_SB2_n715) );
  NAND3_X1 R2_SB_SB2_U426 ( .A1(R2_SB_SB2_n717), .A2(R2_SB_SB2_n716), .A3(
        R2_SB_SB2_n715), .ZN(R2_SB_SB2_n737) );
  NAND4_X1 R2_SB_SB2_U425 ( .A1(R2_SB_SB2_n741), .A2(R2_SB_SB2_n740), .A3(
        R2_SB_SB2_n739), .A4(R2_SB_SB2_n738), .ZN(R2_SB_n319) );
  NAND3_X1 R2_SB_SB2_U424 ( .A1(R2_SB_n328), .A2(R2_SB_SB2_n854), .A3(
        R2_SB_SB2_n795), .ZN(R2_SB_SB2_n762) );
  NAND3_X1 R2_SB_SB2_U423 ( .A1(R2_SB_SB2_n763), .A2(R2_SB_SB2_n762), .A3(
        R2_SB_SB2_n761), .ZN(R2_SB_SB2_n764) );
  NAND3_X1 R2_SB_SB2_U422 ( .A1(R2_SB_n327), .A2(R2_SB_SB2_n854), .A3(
        R2_SB_SB2_n771), .ZN(R2_SB_SB2_n777) );
  NAND3_X1 R2_SB_SB2_U421 ( .A1(R2_SB_SB2_n817), .A2(R2_SB_SB2_n816), .A3(
        R2_SB_SB2_n815), .ZN(R2_SB_SB2_n820) );
  NAND4_X1 R2_SB_SB2_U420 ( .A1(R2_SB_SB2_n825), .A2(R2_SB_SB2_n824), .A3(
        R2_SB_SB2_n823), .A4(R2_SB_SB2_n822), .ZN(R2_SB_n320) );
  NOR2_X2 R2_SB_SB2_U264 ( .A1(R2_SB_SB2_n830), .A2(R2_SB_SB2_n843), .ZN(
        R2_SB_SB2_n758) );
  INV_X1 R2_SB_SB3_U466 ( .A(R2_SB_SB3_n453), .ZN(R2_SB_SB3_n452) );
  INV_X1 R2_SB_SB3_U465 ( .A(R2_SB_n306), .ZN(R2_SB_SB3_n89) );
  INV_X1 R2_SB_SB3_U419 ( .A(R2_SB_n305), .ZN(R2_SB_SB3_n453) );
  NAND2_X1 R2_SB_SB3_U418 ( .A1(R2_SB_n306), .A2(R2_SB_n311), .ZN(
        R2_SB_SB3_n705) );
  AOI22_X1 R2_SB_SB3_U417 ( .A1(R2_SB_SB3_n779), .A2(R2_SB_SB3_n760), .B1(
        R2_SB_SB3_n877), .B2(R2_SB_SB3_n792), .ZN(R2_SB_SB3_n761) );
  OAI21_X1 R2_SB_SB3_U416 ( .B1(R2_SB_SB3_n759), .B2(R2_SB_SB3_n900), .A(
        R2_SB_SB3_n758), .ZN(R2_SB_SB3_n763) );
  AOI222_X1 R2_SB_SB3_U415 ( .A1(R2_SB_SB3_n742), .A2(R2_SB_n310), .B1(
        R2_SB_SB3_n778), .B2(R2_SB_SB3_n748), .C1(R2_SB_SB3_n747), .C2(
        R2_SB_SB3_n656), .ZN(R2_SB_SB3_n657) );
  NAND2_X1 R2_SB_SB3_U414 ( .A1(R2_SB_SB3_n743), .A2(R2_SB_n312), .ZN(
        R2_SB_SB3_n472) );
  AOI21_X1 R2_SB_SB3_U413 ( .B1(R2_SB_SB3_n835), .B2(R2_SB_SB3_n837), .A(
        R2_SB_SB3_n859), .ZN(R2_SB_SB3_n474) );
  OAI21_X1 R2_SB_SB3_U412 ( .B1(R2_SB_SB3_n474), .B2(R2_SB_SB3_n473), .A(
        R2_SB_SB3_n813), .ZN(R2_SB_SB3_n475) );
  OAI22_X1 R2_SB_SB3_U411 ( .A1(R2_SB_SB3_n829), .A2(R2_SB_SB3_n847), .B1(
        R2_SB_SB3_n845), .B2(R2_SB_SB3_n826), .ZN(R2_SB_SB3_n714) );
  NOR2_X1 R2_SB_SB3_U410 ( .A1(R2_SB_n312), .A2(R2_SB_SB3_n863), .ZN(
        R2_SB_SB3_n535) );
  OAI21_X1 R2_SB_SB3_U409 ( .B1(R2_SB_SB3_n855), .B2(R2_SB_SB3_n829), .A(
        R2_SB_SB3_n745), .ZN(R2_SB_SB3_n746) );
  AOI221_X1 R2_SB_SB3_U408 ( .B1(R2_SB_SB3_n805), .B2(R2_SB_SB3_n748), .C1(
        R2_SB_SB3_n747), .C2(R2_SB_SB3_n780), .A(R2_SB_SB3_n746), .ZN(
        R2_SB_SB3_n749) );
  AOI22_X1 R2_SB_SB3_U407 ( .A1(R2_SB_SB3_n742), .A2(R2_SB_n310), .B1(
        R2_SB_SB3_n778), .B2(R2_SB_SB3_n771), .ZN(R2_SB_SB3_n750) );
  OAI211_X1 R2_SB_SB3_U406 ( .C1(R2_SB_SB3_n828), .C2(R2_SB_SB3_n847), .A(
        R2_SB_SB3_n750), .B(R2_SB_SB3_n749), .ZN(R2_SB_SB3_n751) );
  NOR2_X1 R2_SB_SB3_U405 ( .A1(R2_SB_n310), .A2(R2_SB_SB3_n830), .ZN(
        R2_SB_SB3_n724) );
  NOR2_X1 R2_SB_SB3_U404 ( .A1(R2_SB_SB3_n826), .A2(R2_SB_n308), .ZN(
        R2_SB_SB3_n463) );
  OAI22_X1 R2_SB_SB3_U403 ( .A1(R2_SB_n312), .A2(R2_SB_SB3_n876), .B1(
        R2_SB_SB3_n858), .B2(R2_SB_SB3_n901), .ZN(R2_SB_SB3_n760) );
  NOR3_X1 R2_SB_SB3_U402 ( .A1(R2_SB_SB3_n890), .A2(R2_SB_n310), .A3(
        R2_SB_n306), .ZN(R2_SB_SB3_n613) );
  OAI22_X1 R2_SB_SB3_U401 ( .A1(R2_SB_SB3_n89), .A2(R2_SB_SB3_n898), .B1(
        R2_SB_SB3_n628), .B2(R2_SB_SB3_n907), .ZN(R2_SB_SB3_n614) );
  NOR3_X1 R2_SB_SB3_U400 ( .A1(R2_SB_SB3_n614), .A2(R2_SB_SB3_n722), .A3(
        R2_SB_SB3_n613), .ZN(R2_SB_SB3_n623) );
  NOR3_X1 R2_SB_SB3_U399 ( .A1(R2_SB_SB3_n863), .A2(R2_SB_n312), .A3(
        R2_SB_SB3_n814), .ZN(R2_SB_SB3_n797) );
  AOI22_X1 R2_SB_SB3_U398 ( .A1(R2_SB_SB3_n628), .A2(R2_SB_SB3_n627), .B1(
        R2_SB_n307), .B2(R2_SB_SB3_n730), .ZN(R2_SB_SB3_n630) );
  OAI222_X1 R2_SB_SB3_U397 ( .A1(R2_SB_SB3_n837), .A2(R2_SB_SB3_n573), .B1(
        R2_SB_n305), .B2(R2_SB_SB3_n468), .C1(R2_SB_n306), .C2(R2_SB_SB3_n677), 
        .ZN(R2_SB_SB3_n483) );
  OAI221_X1 R2_SB_SB3_U396 ( .B1(R2_SB_n308), .B2(R2_SB_SB3_n581), .C1(
        R2_SB_SB3_n476), .C2(R2_SB_SB3_n878), .A(R2_SB_SB3_n475), .ZN(
        R2_SB_SB3_n482) );
  OAI22_X1 R2_SB_SB3_U395 ( .A1(R2_SB_SB3_n840), .A2(R2_SB_SB3_n800), .B1(
        R2_SB_SB3_n480), .B2(R2_SB_SB3_n453), .ZN(R2_SB_SB3_n481) );
  NOR4_X1 R2_SB_SB3_U394 ( .A1(R2_SB_SB3_n484), .A2(R2_SB_SB3_n483), .A3(
        R2_SB_SB3_n482), .A4(R2_SB_SB3_n481), .ZN(R2_SB_SB3_n485) );
  NOR2_X1 R2_SB_SB3_U393 ( .A1(R2_SB_SB3_n868), .A2(R2_SB_n312), .ZN(
        R2_SB_SB3_n680) );
  NOR2_X1 R2_SB_SB3_U392 ( .A1(R2_SB_n307), .A2(R2_SB_n309), .ZN(
        R2_SB_SB3_n646) );
  NAND2_X1 R2_SB_SB3_U391 ( .A1(R2_SB_n310), .A2(R2_SB_SB3_n872), .ZN(
        R2_SB_SB3_n770) );
  NOR2_X1 R2_SB_SB3_U390 ( .A1(R2_SB_SB3_n895), .A2(R2_SB_n308), .ZN(
        R2_SB_SB3_n783) );
  NOR2_X1 R2_SB_SB3_U389 ( .A1(R2_SB_n309), .A2(R2_SB_n310), .ZN(
        R2_SB_SB3_n617) );
  NOR2_X1 R2_SB_SB3_U388 ( .A1(R2_SB_SB3_n854), .A2(R2_SB_n307), .ZN(
        R2_SB_SB3_n811) );
  INV_X1 R2_SB_SB3_U387 ( .A(R2_SB_n312), .ZN(R2_SB_SB3_n881) );
  AOI22_X1 R2_SB_SB3_U386 ( .A1(R2_SB_n307), .A2(R2_SB_SB3_n638), .B1(
        R2_SB_SB3_n795), .B2(R2_SB_SB3_n713), .ZN(R2_SB_SB3_n711) );
  NOR2_X1 R2_SB_SB3_U385 ( .A1(R2_SB_SB3_n854), .A2(R2_SB_n310), .ZN(
        R2_SB_SB3_n694) );
  NAND2_X1 R2_SB_SB3_U384 ( .A1(R2_SB_n307), .A2(R2_SB_n310), .ZN(
        R2_SB_SB3_n608) );
  OAI221_X1 R2_SB_SB3_U383 ( .B1(R2_SB_n307), .B2(R2_SB_SB3_n551), .C1(
        R2_SB_SB3_n550), .C2(R2_SB_SB3_n910), .A(R2_SB_SB3_n902), .ZN(
        R2_SB_SB3_n552) );
  OAI221_X1 R2_SB_SB3_U382 ( .B1(R2_SB_SB3_n864), .B2(R2_SB_SB3_n838), .C1(
        R2_SB_SB3_n827), .C2(R2_SB_SB3_n849), .A(R2_SB_SB3_n615), .ZN(
        R2_SB_SB3_n553) );
  OAI221_X1 R2_SB_SB3_U381 ( .B1(R2_SB_SB3_n864), .B2(R2_SB_SB3_n835), .C1(
        R2_SB_SB3_n832), .C2(R2_SB_SB3_n853), .A(R2_SB_SB3_n546), .ZN(
        R2_SB_SB3_n554) );
  AOI221_X1 R2_SB_SB3_U380 ( .B1(R2_SB_SB3_n752), .B2(R2_SB_SB3_n554), .C1(
        R2_SB_SB3_n702), .C2(R2_SB_SB3_n553), .A(R2_SB_SB3_n552), .ZN(
        R2_SB_SB3_n559) );
  OAI22_X1 R2_SB_SB3_U379 ( .A1(R2_SB_SB3_n583), .A2(R2_SB_SB3_n826), .B1(
        R2_SB_SB3_n838), .B2(R2_SB_SB3_n891), .ZN(R2_SB_SB3_n584) );
  OAI211_X1 R2_SB_SB3_U378 ( .C1(R2_SB_SB3_n453), .C2(R2_SB_SB3_n844), .A(
        R2_SB_SB3_n835), .B(R2_SB_SB3_n847), .ZN(R2_SB_SB3_n585) );
  OAI211_X1 R2_SB_SB3_U377 ( .C1(R2_SB_n305), .C2(R2_SB_SB3_n898), .A(
        R2_SB_SB3_n582), .B(R2_SB_SB3_n581), .ZN(R2_SB_SB3_n586) );
  AOI221_X1 R2_SB_SB3_U376 ( .B1(R2_SB_n307), .B2(R2_SB_SB3_n586), .C1(
        R2_SB_SB3_n755), .C2(R2_SB_SB3_n585), .A(R2_SB_SB3_n584), .ZN(
        R2_SB_SB3_n599) );
  OAI221_X1 R2_SB_SB3_U375 ( .B1(R2_SB_SB3_n840), .B2(R2_SB_SB3_n859), .C1(
        R2_SB_SB3_n863), .C2(R2_SB_SB3_n834), .A(R2_SB_SB3_n574), .ZN(
        R2_SB_SB3_n580) );
  OAI22_X1 R2_SB_SB3_U374 ( .A1(R2_SB_n308), .A2(R2_SB_SB3_n578), .B1(
        R2_SB_SB3_n577), .B2(R2_SB_SB3_n831), .ZN(R2_SB_SB3_n579) );
  INV_X1 R2_SB_SB3_U373 ( .A(R2_SB_SB3_n573), .ZN(R2_SB_SB3_n889) );
  AOI221_X1 R2_SB_SB3_U372 ( .B1(R2_SB_SB3_n889), .B2(R2_SB_SB3_n696), .C1(
        R2_SB_SB3_n752), .C2(R2_SB_SB3_n580), .A(R2_SB_SB3_n579), .ZN(
        R2_SB_SB3_n600) );
  NOR2_X1 R2_SB_SB3_U371 ( .A1(R2_SB_n308), .A2(R2_SB_n309), .ZN(
        R2_SB_SB3_n656) );
  INV_X1 R2_SB_SB3_U370 ( .A(R2_SB_n311), .ZN(R2_SB_SB3_n872) );
  NOR3_X1 R2_SB_SB3_U369 ( .A1(R2_SB_SB3_n850), .A2(R2_SB_n309), .A3(
        R2_SB_SB3_n881), .ZN(R2_SB_SB3_n556) );
  NOR2_X1 R2_SB_SB3_U368 ( .A1(R2_SB_SB3_n830), .A2(R2_SB_n309), .ZN(
        R2_SB_SB3_n678) );
  AOI221_X1 R2_SB_SB3_U367 ( .B1(R2_SB_SB3_n806), .B2(R2_SB_SB3_n89), .C1(
        R2_SB_SB3_n805), .C2(R2_SB_SB3_n804), .A(R2_SB_SB3_n803), .ZN(
        R2_SB_SB3_n807) );
  AOI211_X1 R2_SB_SB3_U366 ( .C1(R2_SB_SB3_n799), .C2(R2_SB_SB3_n798), .A(
        R2_SB_SB3_n797), .B(R2_SB_SB3_n796), .ZN(R2_SB_SB3_n808) );
  AOI22_X1 R2_SB_SB3_U365 ( .A1(R2_SB_SB3_n793), .A2(R2_SB_SB3_n792), .B1(
        R2_SB_SB3_n791), .B2(R2_SB_SB3_n790), .ZN(R2_SB_SB3_n809) );
  OAI221_X1 R2_SB_SB3_U364 ( .B1(R2_SB_n311), .B2(R2_SB_SB3_n809), .C1(
        R2_SB_SB3_n808), .C2(R2_SB_SB3_n859), .A(R2_SB_SB3_n807), .ZN(
        R2_SB_SB3_n821) );
  NOR2_X1 R2_SB_SB3_U363 ( .A1(R2_SB_n312), .A2(R2_SB_n309), .ZN(
        R2_SB_SB3_n489) );
  OAI21_X1 R2_SB_SB3_U362 ( .B1(R2_SB_SB3_n864), .B2(R2_SB_SB3_n878), .A(
        R2_SB_SB3_n894), .ZN(R2_SB_SB3_n490) );
  AOI221_X1 R2_SB_SB3_U361 ( .B1(R2_SB_SB3_n779), .B2(R2_SB_SB3_n490), .C1(
        R2_SB_SB3_n489), .C2(R2_SB_SB3_n782), .A(R2_SB_SB3_n756), .ZN(
        R2_SB_SB3_n491) );
  AOI222_X1 R2_SB_SB3_U360 ( .A1(R2_SB_SB3_n789), .A2(R2_SB_SB3_n772), .B1(
        R2_SB_SB3_n646), .B2(R2_SB_SB3_n813), .C1(R2_SB_SB3_n709), .C2(
        R2_SB_SB3_n811), .ZN(R2_SB_SB3_n647) );
  OAI221_X1 R2_SB_SB3_U359 ( .B1(R2_SB_n306), .B2(R2_SB_SB3_n884), .C1(
        R2_SB_SB3_n453), .C2(R2_SB_SB3_n880), .A(R2_SB_SB3_n649), .ZN(
        R2_SB_SB3_n650) );
  OAI221_X1 R2_SB_SB3_U358 ( .B1(R2_SB_n308), .B2(R2_SB_SB3_n648), .C1(
        R2_SB_SB3_n845), .C2(R2_SB_SB3_n868), .A(R2_SB_SB3_n647), .ZN(
        R2_SB_SB3_n652) );
  AOI222_X1 R2_SB_SB3_U357 ( .A1(R2_SB_SB3_n781), .A2(R2_SB_SB3_n652), .B1(
        R2_SB_SB3_n651), .B2(R2_SB_SB3_n730), .C1(R2_SB_SB3_n782), .C2(
        R2_SB_SB3_n650), .ZN(R2_SB_SB3_n693) );
  NOR2_X1 R2_SB_SB3_U356 ( .A1(R2_SB_SB3_n863), .A2(R2_SB_n308), .ZN(
        R2_SB_SB3_n618) );
  NOR3_X1 R2_SB_SB3_U355 ( .A1(R2_SB_SB3_n840), .A2(R2_SB_n311), .A3(
        R2_SB_SB3_n869), .ZN(R2_SB_SB3_n575) );
  AOI221_X1 R2_SB_SB3_U354 ( .B1(R2_SB_SB3_n591), .B2(R2_SB_SB3_n453), .C1(
        R2_SB_SB3_n576), .C2(R2_SB_SB3_n684), .A(R2_SB_SB3_n575), .ZN(
        R2_SB_SB3_n578) );
  OAI211_X1 R2_SB_SB3_U353 ( .C1(R2_SB_n310), .C2(R2_SB_SB3_n848), .A(
        R2_SB_SB3_n860), .B(R2_SB_SB3_n853), .ZN(R2_SB_SB3_n662) );
  OAI21_X1 R2_SB_SB3_U352 ( .B1(R2_SB_SB3_n876), .B2(R2_SB_SB3_n853), .A(
        R2_SB_SB3_n908), .ZN(R2_SB_SB3_n663) );
  AOI221_X1 R2_SB_SB3_U351 ( .B1(R2_SB_SB3_n779), .B2(R2_SB_SB3_n663), .C1(
        R2_SB_SB3_n702), .C2(R2_SB_SB3_n662), .A(R2_SB_SB3_n661), .ZN(
        R2_SB_SB3_n664) );
  OAI222_X1 R2_SB_SB3_U350 ( .A1(R2_SB_SB3_n718), .A2(R2_SB_SB3_n907), .B1(
        R2_SB_SB3_n452), .B2(R2_SB_SB3_n664), .C1(R2_SB_SB3_n832), .C2(
        R2_SB_SB3_n802), .ZN(R2_SB_SB3_n667) );
  NOR3_X1 R2_SB_SB3_U349 ( .A1(R2_SB_SB3_n849), .A2(R2_SB_n312), .A3(
        R2_SB_SB3_n854), .ZN(R2_SB_SB3_n605) );
  OAI22_X1 R2_SB_SB3_U348 ( .A1(R2_SB_n311), .A2(R2_SB_n309), .B1(R2_SB_n310), 
        .B2(R2_SB_SB3_n883), .ZN(R2_SB_SB3_n606) );
  AOI221_X1 R2_SB_SB3_U347 ( .B1(R2_SB_SB3_n755), .B2(R2_SB_SB3_n791), .C1(
        R2_SB_SB3_n758), .C2(R2_SB_SB3_n606), .A(R2_SB_SB3_n605), .ZN(
        R2_SB_SB3_n607) );
  NOR2_X1 R2_SB_SB3_U346 ( .A1(R2_SB_SB3_n452), .A2(R2_SB_n307), .ZN(
        R2_SB_SB3_n794) );
  NOR2_X1 R2_SB_SB3_U345 ( .A1(R2_SB_n310), .A2(R2_SB_n312), .ZN(
        R2_SB_SB3_n709) );
  NOR2_X1 R2_SB_SB3_U344 ( .A1(R2_SB_SB3_n830), .A2(R2_SB_n308), .ZN(
        R2_SB_SB3_n782) );
  NOR3_X1 R2_SB_SB3_U343 ( .A1(R2_SB_SB3_n901), .A2(R2_SB_n311), .A3(
        R2_SB_SB3_n843), .ZN(R2_SB_SB3_n729) );
  AOI221_X1 R2_SB_SB3_U342 ( .B1(R2_SB_SB3_n805), .B2(R2_SB_SB3_n813), .C1(
        R2_SB_SB3_n789), .C2(R2_SB_SB3_n728), .A(R2_SB_SB3_n727), .ZN(
        R2_SB_SB3_n732) );
  AOI211_X1 R2_SB_SB3_U341 ( .C1(R2_SB_SB3_n752), .C2(R2_SB_SB3_n730), .A(
        R2_SB_SB3_n759), .B(R2_SB_SB3_n729), .ZN(R2_SB_SB3_n731) );
  OAI222_X1 R2_SB_SB3_U340 ( .A1(R2_SB_SB3_n733), .A2(R2_SB_SB3_n839), .B1(
        R2_SB_SB3_n732), .B2(R2_SB_SB3_n837), .C1(R2_SB_SB3_n731), .C2(
        R2_SB_SB3_n835), .ZN(R2_SB_SB3_n734) );
  NOR2_X1 R2_SB_SB3_U339 ( .A1(R2_SB_SB3_n854), .A2(R2_SB_n308), .ZN(
        R2_SB_SB3_n805) );
  NOR2_X1 R2_SB_SB3_U338 ( .A1(R2_SB_SB3_n872), .A2(R2_SB_n310), .ZN(
        R2_SB_SB3_n767) );
  INV_X1 R2_SB_SB3_U337 ( .A(R2_SB_n307), .ZN(R2_SB_SB3_n830) );
  NOR2_X1 R2_SB_SB3_U336 ( .A1(R2_SB_n311), .A2(R2_SB_n312), .ZN(
        R2_SB_SB3_n702) );
  NOR2_X1 R2_SB_SB3_U335 ( .A1(R2_SB_n306), .A2(R2_SB_n307), .ZN(
        R2_SB_SB3_n795) );
  NOR2_X1 R2_SB_SB3_U334 ( .A1(R2_SB_n310), .A2(R2_SB_n311), .ZN(
        R2_SB_SB3_n813) );
  NOR3_X1 R2_SB_SB3_U333 ( .A1(R2_SB_SB3_n833), .A2(R2_SB_n308), .A3(
        R2_SB_SB3_n885), .ZN(R2_SB_SB3_n639) );
  INV_X1 R2_SB_SB3_U332 ( .A(R2_SB_n309), .ZN(R2_SB_SB3_n854) );
  NOR2_X1 R2_SB_SB3_U331 ( .A1(R2_SB_SB3_n843), .A2(R2_SB_n307), .ZN(
        R2_SB_SB3_n792) );
  INV_X1 R2_SB_SB3_U330 ( .A(R2_SB_n310), .ZN(R2_SB_SB3_n863) );
  NAND2_X1 R2_SB_SB3_U329 ( .A1(R2_SB_SB3_n791), .A2(R2_SB_SB3_n772), .ZN(
        R2_SB_SB3_n775) );
  OAI21_X1 R2_SB_SB3_U328 ( .B1(R2_SB_SB3_n775), .B2(R2_SB_SB3_n774), .A(
        R2_SB_SB3_n773), .ZN(R2_SB_SB3_n776) );
  INV_X1 R2_SB_SB3_U327 ( .A(R2_SB_SB3_n776), .ZN(R2_SB_SB3_n887) );
  INV_X1 R2_SB_SB3_U326 ( .A(R2_SB_SB3_n783), .ZN(R2_SB_SB3_n897) );
  INV_X1 R2_SB_SB3_U325 ( .A(R2_SB_SB3_n678), .ZN(R2_SB_SB3_n860) );
  INV_X1 R2_SB_SB3_U324 ( .A(R2_SB_SB3_n811), .ZN(R2_SB_SB3_n855) );
  INV_X1 R2_SB_SB3_U323 ( .A(R2_SB_SB3_n463), .ZN(R2_SB_SB3_n842) );
  INV_X1 R2_SB_SB3_U322 ( .A(R2_SB_SB3_n711), .ZN(R2_SB_SB3_n909) );
  NAND2_X1 R2_SB_SB3_U321 ( .A1(R2_SB_SB3_n678), .A2(R2_SB_SB3_n781), .ZN(
        R2_SB_SB3_n615) );
  NAND2_X1 R2_SB_SB3_U320 ( .A1(R2_SB_SB3_n680), .A2(R2_SB_SB3_n810), .ZN(
        R2_SB_SB3_n581) );
  NAND2_X1 R2_SB_SB3_U319 ( .A1(R2_SB_SB3_n772), .A2(R2_SB_SB3_n684), .ZN(
        R2_SB_SB3_n785) );
  NAND2_X1 R2_SB_SB3_U318 ( .A1(R2_SB_SB3_n670), .A2(R2_SB_SB3_n881), .ZN(
        R2_SB_SB3_n773) );
  NAND2_X1 R2_SB_SB3_U317 ( .A1(R2_SB_SB3_n670), .A2(R2_SB_SB3_n872), .ZN(
        R2_SB_SB3_n801) );
  NAND2_X1 R2_SB_SB3_U316 ( .A1(R2_SB_SB3_n452), .A2(R2_SB_SB3_n843), .ZN(
        R2_SB_SB3_n548) );
  NOR2_X1 R2_SB_SB3_U315 ( .A1(R2_SB_SB3_n854), .A2(R2_SB_SB3_n827), .ZN(
        R2_SB_SB3_n793) );
  OAI21_X1 R2_SB_SB3_U314 ( .B1(R2_SB_SB3_n718), .B2(R2_SB_SB3_n588), .A(
        R2_SB_SB3_n587), .ZN(R2_SB_SB3_n597) );
  AOI22_X1 R2_SB_SB3_U313 ( .A1(R2_SB_SB3_n753), .A2(R2_SB_SB3_n771), .B1(
        R2_SB_SB3_n752), .B2(R2_SB_SB3_n751), .ZN(R2_SB_SB3_n825) );
  AOI22_X1 R2_SB_SB3_U312 ( .A1(R2_SB_n306), .A2(R2_SB_SB3_n765), .B1(
        R2_SB_SB3_n764), .B2(R2_SB_SB3_n453), .ZN(R2_SB_SB3_n824) );
  NOR4_X1 R2_SB_SB3_U311 ( .A1(R2_SB_SB3_n464), .A2(R2_SB_SB3_n886), .A3(
        R2_SB_SB3_n555), .A4(R2_SB_SB3_n639), .ZN(R2_SB_SB3_n486) );
  AOI211_X1 R2_SB_SB3_U310 ( .C1(R2_SB_SB3_n684), .C2(R2_SB_SB3_n462), .A(
        R2_SB_SB3_n461), .B(R2_SB_SB3_n460), .ZN(R2_SB_SB3_n487) );
  AOI221_X1 R2_SB_SB3_U309 ( .B1(R2_SB_SB3_n810), .B2(R2_SB_SB3_n533), .C1(
        R2_SB_SB3_n565), .C2(R2_SB_n306), .A(R2_SB_SB3_n532), .ZN(
        R2_SB_SB3_n561) );
  NOR4_X1 R2_SB_SB3_U308 ( .A1(R2_SB_SB3_n557), .A2(R2_SB_SB3_n556), .A3(
        R2_SB_SB3_n555), .A4(R2_SB_SB3_n674), .ZN(R2_SB_SB3_n558) );
  AOI221_X1 R2_SB_SB3_U307 ( .B1(R2_SB_SB3_n772), .B2(R2_SB_SB3_n572), .C1(
        R2_SB_SB3_n753), .C2(R2_SB_SB3_n758), .A(R2_SB_SB3_n571), .ZN(
        R2_SB_SB3_n601) );
  AOI211_X1 R2_SB_SB3_U306 ( .C1(R2_SB_SB3_n597), .C2(R2_SB_SB3_n453), .A(
        R2_SB_SB3_n596), .B(R2_SB_SB3_n595), .ZN(R2_SB_SB3_n598) );
  AOI221_X1 R2_SB_SB3_U305 ( .B1(R2_SB_SB3_n604), .B2(R2_SB_SB3_n877), .C1(
        R2_SB_SB3_n603), .C2(R2_SB_SB3_n679), .A(R2_SB_SB3_n602), .ZN(
        R2_SB_SB3_n645) );
  NOR4_X1 R2_SB_SB3_U304 ( .A1(R2_SB_SB3_n641), .A2(R2_SB_SB3_n640), .A3(
        R2_SB_SB3_n639), .A4(R2_SB_SB3_n673), .ZN(R2_SB_SB3_n642) );
  OAI21_X1 R2_SB_SB3_U303 ( .B1(R2_SB_SB3_n810), .B2(R2_SB_SB3_n744), .A(
        R2_SB_SB3_n743), .ZN(R2_SB_SB3_n745) );
  NOR4_X1 R2_SB_SB3_U302 ( .A1(R2_SB_SB3_n737), .A2(R2_SB_SB3_n736), .A3(
        R2_SB_SB3_n735), .A4(R2_SB_SB3_n734), .ZN(R2_SB_SB3_n738) );
  AOI211_X1 R2_SB_SB3_U301 ( .C1(R2_SB_SB3_n713), .C2(R2_SB_SB3_n758), .A(
        R2_SB_SB3_n712), .B(R2_SB_SB3_n909), .ZN(R2_SB_SB3_n739) );
  NOR4_X1 R2_SB_SB3_U300 ( .A1(R2_SB_SB3_n689), .A2(R2_SB_SB3_n688), .A3(
        R2_SB_SB3_n687), .A4(R2_SB_SB3_n686), .ZN(R2_SB_SB3_n690) );
  AOI211_X1 R2_SB_SB3_U299 ( .C1(R2_SB_SB3_n752), .C2(R2_SB_SB3_n668), .A(
        R2_SB_SB3_n667), .B(R2_SB_SB3_n666), .ZN(R2_SB_SB3_n691) );
  AOI221_X1 R2_SB_SB3_U298 ( .B1(R2_SB_SB3_n565), .B2(R2_SB_SB3_n766), .C1(
        R2_SB_SB3_n759), .C2(R2_SB_SB3_n791), .A(R2_SB_SB3_n513), .ZN(
        R2_SB_SB3_n525) );
  NOR4_X1 R2_SB_SB3_U297 ( .A1(R2_SB_SB3_n523), .A2(R2_SB_SB3_n522), .A3(
        R2_SB_SB3_n521), .A4(R2_SB_SB3_n520), .ZN(R2_SB_SB3_n524) );
  OAI221_X1 R2_SB_SB3_U296 ( .B1(R2_SB_SB3_n849), .B2(R2_SB_SB3_n770), .C1(
        R2_SB_SB3_n883), .C2(R2_SB_SB3_n608), .A(R2_SB_SB3_n567), .ZN(
        R2_SB_SB3_n568) );
  OAI21_X1 R2_SB_SB3_U295 ( .B1(R2_SB_SB3_n569), .B2(R2_SB_SB3_n568), .A(
        R2_SB_SB3_n781), .ZN(R2_SB_SB3_n570) );
  OAI21_X1 R2_SB_SB3_U294 ( .B1(R2_SB_SB3_n839), .B2(R2_SB_SB3_n892), .A(
        R2_SB_SB3_n570), .ZN(R2_SB_SB3_n571) );
  INV_X1 R2_SB_SB3_U293 ( .A(R2_SB_SB3_n780), .ZN(R2_SB_SB3_n870) );
  OAI21_X1 R2_SB_SB3_U292 ( .B1(R2_SB_SB3_n778), .B2(R2_SB_SB3_n744), .A(
        R2_SB_SB3_n696), .ZN(R2_SB_SB3_n508) );
  OAI211_X1 R2_SB_SB3_U291 ( .C1(R2_SB_SB3_n813), .C2(R2_SB_SB3_n812), .A(
        R2_SB_SB3_n811), .B(R2_SB_SB3_n810), .ZN(R2_SB_SB3_n817) );
  INV_X1 R2_SB_SB3_U290 ( .A(R2_SB_SB3_n743), .ZN(R2_SB_SB3_n851) );
  AND3_X1 R2_SB_SB3_U289 ( .A1(R2_SB_SB3_n779), .A2(R2_SB_SB3_n812), .A3(
        R2_SB_SB3_n656), .ZN(R2_SB_SB3_n87) );
  NOR3_X1 R2_SB_SB3_U288 ( .A1(R2_SB_SB3_n858), .A2(R2_SB_SB3_n665), .A3(
        R2_SB_SB3_n890), .ZN(R2_SB_SB3_n13) );
  OR3_X1 R2_SB_SB3_U287 ( .A1(R2_SB_SB3_n13), .A2(R2_SB_SB3_n675), .A3(
        R2_SB_SB3_n87), .ZN(R2_SB_SB3_n464) );
  OAI22_X1 R2_SB_SB3_U286 ( .A1(R2_SB_SB3_n872), .A2(R2_SB_SB3_n857), .B1(
        R2_SB_SB3_n854), .B2(R2_SB_SB3_n876), .ZN(R2_SB_SB3_n547) );
  INV_X1 R2_SB_SB3_U285 ( .A(R2_SB_SB3_n582), .ZN(R2_SB_SB3_n911) );
  AOI21_X1 R2_SB_SB3_U284 ( .B1(R2_SB_SB3_n781), .B2(R2_SB_SB3_n547), .A(
        R2_SB_SB3_n911), .ZN(R2_SB_SB3_n551) );
  AOI21_X1 R2_SB_SB3_U283 ( .B1(R2_SB_SB3_n754), .B2(R2_SB_SB3_n758), .A(
        R2_SB_SB3_n467), .ZN(R2_SB_SB3_n468) );
  AOI21_X1 R2_SB_SB3_U282 ( .B1(R2_SB_SB3_n778), .B2(R2_SB_SB3_n453), .A(
        R2_SB_SB3_n789), .ZN(R2_SB_SB3_n700) );
  AOI22_X1 R2_SB_SB3_U281 ( .A1(R2_SB_SB3_n725), .A2(R2_SB_SB3_n617), .B1(
        R2_SB_SB3_n766), .B2(R2_SB_SB3_n730), .ZN(R2_SB_SB3_n562) );
  AOI21_X1 R2_SB_SB3_U280 ( .B1(R2_SB_SB3_n743), .B2(R2_SB_n306), .A(
        R2_SB_SB3_n747), .ZN(R2_SB_SB3_n564) );
  OAI21_X1 R2_SB_SB3_U279 ( .B1(R2_SB_SB3_n684), .B2(R2_SB_SB3_n799), .A(
        R2_SB_SB3_n780), .ZN(R2_SB_SB3_n563) );
  OAI211_X1 R2_SB_SB3_U278 ( .C1(R2_SB_SB3_n564), .C2(R2_SB_SB3_n868), .A(
        R2_SB_SB3_n563), .B(R2_SB_SB3_n562), .ZN(R2_SB_SB3_n572) );
  OAI21_X1 R2_SB_SB3_U277 ( .B1(R2_SB_SB3_n905), .B2(R2_SB_SB3_n859), .A(
        R2_SB_SB3_n895), .ZN(R2_SB_SB3_n529) );
  AOI211_X1 R2_SB_SB3_U276 ( .C1(R2_SB_SB3_n529), .C2(R2_SB_SB3_n830), .A(
        R2_SB_SB3_n633), .B(R2_SB_SB3_n528), .ZN(R2_SB_SB3_n530) );
  AOI22_X1 R2_SB_SB3_U275 ( .A1(R2_SB_SB3_n680), .A2(R2_SB_SB3_n843), .B1(
        R2_SB_SB3_n678), .B2(R2_SB_SB3_n772), .ZN(R2_SB_SB3_n531) );
  OAI211_X1 R2_SB_SB3_U274 ( .C1(R2_SB_SB3_n905), .C2(R2_SB_SB3_n864), .A(
        R2_SB_SB3_n531), .B(R2_SB_SB3_n530), .ZN(R2_SB_SB3_n533) );
  OAI21_X1 R2_SB_SB3_U273 ( .B1(R2_SB_SB3_n755), .B2(R2_SB_SB3_n754), .A(
        R2_SB_SB3_n782), .ZN(R2_SB_SB3_n757) );
  INV_X1 R2_SB_SB3_U272 ( .A(R2_SB_SB3_n756), .ZN(R2_SB_SB3_n899) );
  OAI211_X1 R2_SB_SB3_U271 ( .C1(R2_SB_SB3_n845), .C2(R2_SB_SB3_n880), .A(
        R2_SB_SB3_n757), .B(R2_SB_SB3_n899), .ZN(R2_SB_SB3_n765) );
  INV_X1 R2_SB_SB3_U270 ( .A(R2_SB_SB3_n696), .ZN(R2_SB_SB3_n836) );
  AOI21_X1 R2_SB_SB3_U269 ( .B1(R2_SB_SB3_n843), .B2(R2_SB_SB3_n835), .A(
        R2_SB_SB3_n879), .ZN(R2_SB_SB3_n595) );
  NAND2_X1 R2_SB_SB3_U268 ( .A1(R2_SB_SB3_n634), .A2(R2_SB_SB3_n805), .ZN(
        R2_SB_SB3_n800) );
  NAND2_X1 R2_SB_SB3_U267 ( .A1(R2_SB_SB3_n772), .A2(R2_SB_SB3_n507), .ZN(
        R2_SB_SB3_n648) );
  AOI21_X1 R2_SB_SB3_U266 ( .B1(R2_SB_SB3_n849), .B2(R2_SB_SB3_n608), .A(
        R2_SB_SB3_n878), .ZN(R2_SB_SB3_n528) );
  INV_X1 R2_SB_SB3_U265 ( .A(R2_SB_SB3_n794), .ZN(R2_SB_SB3_n837) );
  NOR2_X1 R2_SB_SB3_U263 ( .A1(R2_SB_SB3_n770), .A2(R2_SB_SB3_n833), .ZN(
        R2_SB_SB3_n651) );
  INV_X1 R2_SB_SB3_U262 ( .A(R2_SB_SB3_n798), .ZN(R2_SB_SB3_n901) );
  INV_X1 R2_SB_SB3_U261 ( .A(R2_SB_SB3_n813), .ZN(R2_SB_SB3_n876) );
  AOI22_X1 R2_SB_SB3_U260 ( .A1(R2_SB_SB3_n696), .A2(R2_SB_SB3_n789), .B1(
        R2_SB_SB3_n778), .B2(R2_SB_SB3_n779), .ZN(R2_SB_SB3_n612) );
  AOI22_X1 R2_SB_SB3_U259 ( .A1(R2_SB_SB3_n795), .A2(R2_SB_SB3_n798), .B1(
        R2_SB_SB3_n767), .B2(R2_SB_SB3_n766), .ZN(R2_SB_SB3_n768) );
  NAND2_X1 R2_SB_SB3_U258 ( .A1(R2_SB_SB3_n865), .A2(R2_SB_SB3_n853), .ZN(
        R2_SB_SB3_n495) );
  AOI22_X1 R2_SB_SB3_U257 ( .A1(R2_SB_SB3_n684), .A2(R2_SB_SB3_n495), .B1(
        R2_SB_SB3_n696), .B2(R2_SB_SB3_n618), .ZN(R2_SB_SB3_n496) );
  INV_X1 R2_SB_SB3_U256 ( .A(R2_SB_SB3_n805), .ZN(R2_SB_SB3_n857) );
  NAND2_X1 R2_SB_SB3_U255 ( .A1(R2_SB_SB3_n843), .A2(R2_SB_SB3_n863), .ZN(
        R2_SB_SB3_n774) );
  AOI22_X1 R2_SB_SB3_U254 ( .A1(R2_SB_SB3_n798), .A2(R2_SB_SB3_n627), .B1(
        R2_SB_SB3_n743), .B2(R2_SB_SB3_n752), .ZN(R2_SB_SB3_n567) );
  INV_X1 R2_SB_SB3_U253 ( .A(R2_SB_SB3_n767), .ZN(R2_SB_SB3_n874) );
  NOR2_X1 R2_SB_SB3_U252 ( .A1(R2_SB_SB3_n795), .A2(R2_SB_SB3_n794), .ZN(
        R2_SB_SB3_n814) );
  INV_X1 R2_SB_SB3_U251 ( .A(R2_SB_SB3_n694), .ZN(R2_SB_SB3_n869) );
  NOR2_X1 R2_SB_SB3_U250 ( .A1(R2_SB_SB3_n830), .A2(R2_SB_SB3_n684), .ZN(
        R2_SB_SB3_n665) );
  NOR2_X1 R2_SB_SB3_U249 ( .A1(R2_SB_SB3_n843), .A2(R2_SB_n306), .ZN(
        R2_SB_SB3_n604) );
  NOR2_X1 R2_SB_SB3_U248 ( .A1(R2_SB_SB3_n863), .A2(R2_SB_SB3_n858), .ZN(
        R2_SB_SB3_n790) );
  NAND2_X1 R2_SB_SB3_U247 ( .A1(R2_SB_SB3_n752), .A2(R2_SB_SB3_n507), .ZN(
        R2_SB_SB3_n802) );
  AOI21_X1 R2_SB_SB3_U246 ( .B1(R2_SB_SB3_n789), .B2(R2_SB_SB3_n798), .A(
        R2_SB_SB3_n783), .ZN(R2_SB_SB3_n721) );
  OAI21_X1 R2_SB_SB3_U245 ( .B1(R2_SB_SB3_n747), .B2(R2_SB_SB3_n843), .A(
        R2_SB_SB3_n759), .ZN(R2_SB_SB3_n719) );
  OR3_X1 R2_SB_SB3_U244 ( .A1(R2_SB_SB3_n718), .A2(R2_SB_SB3_n452), .A3(
        R2_SB_SB3_n802), .ZN(R2_SB_SB3_n720) );
  OAI211_X1 R2_SB_SB3_U243 ( .C1(R2_SB_SB3_n721), .C2(R2_SB_SB3_n826), .A(
        R2_SB_SB3_n720), .B(R2_SB_SB3_n719), .ZN(R2_SB_SB3_n736) );
  AOI22_X1 R2_SB_SB3_U242 ( .A1(R2_SB_SB3_n678), .A2(R2_SB_SB3_n767), .B1(
        R2_SB_SB3_n900), .B2(R2_SB_SB3_n843), .ZN(R2_SB_SB3_n683) );
  OAI21_X1 R2_SB_SB3_U241 ( .B1(R2_SB_SB3_n794), .B2(R2_SB_SB3_n791), .A(
        R2_SB_SB3_n882), .ZN(R2_SB_SB3_n681) );
  OAI21_X1 R2_SB_SB3_U240 ( .B1(R2_SB_SB3_n680), .B2(R2_SB_SB3_n679), .A(
        R2_SB_SB3_n696), .ZN(R2_SB_SB3_n682) );
  OAI211_X1 R2_SB_SB3_U239 ( .C1(R2_SB_SB3_n683), .C2(R2_SB_SB3_n829), .A(
        R2_SB_SB3_n682), .B(R2_SB_SB3_n681), .ZN(R2_SB_SB3_n688) );
  NOR3_X1 R2_SB_SB3_U238 ( .A1(R2_SB_SB3_n848), .A2(R2_SB_SB3_n452), .A3(
        R2_SB_SB3_n863), .ZN(R2_SB_SB3_n540) );
  OAI22_X1 R2_SB_SB3_U237 ( .A1(R2_SB_SB3_n858), .A2(R2_SB_SB3_n838), .B1(
        R2_SB_SB3_n857), .B2(R2_SB_SB3_n840), .ZN(R2_SB_SB3_n541) );
  AOI21_X1 R2_SB_SB3_U236 ( .B1(R2_SB_n306), .B2(R2_SB_SB3_n548), .A(
        R2_SB_SB3_n862), .ZN(R2_SB_SB3_n539) );
  NOR3_X1 R2_SB_SB3_U235 ( .A1(R2_SB_SB3_n541), .A2(R2_SB_SB3_n540), .A3(
        R2_SB_SB3_n539), .ZN(R2_SB_SB3_n542) );
  AOI21_X1 R2_SB_SB3_U234 ( .B1(R2_SB_SB3_n730), .B2(R2_SB_SB3_n709), .A(
        R2_SB_SB3_n753), .ZN(R2_SB_SB3_n733) );
  INV_X1 R2_SB_SB3_U233 ( .A(R2_SB_SB3_n791), .ZN(R2_SB_SB3_n840) );
  NOR3_X1 R2_SB_SB3_U232 ( .A1(R2_SB_SB3_n828), .A2(R2_SB_SB3_n856), .A3(
        R2_SB_SB3_n876), .ZN(R2_SB_SB3_n819) );
  AOI21_X1 R2_SB_SB3_U231 ( .B1(R2_SB_SB3_n845), .B2(R2_SB_SB3_n837), .A(
        R2_SB_SB3_n906), .ZN(R2_SB_SB3_n818) );
  NOR4_X1 R2_SB_SB3_U230 ( .A1(R2_SB_SB3_n821), .A2(R2_SB_SB3_n820), .A3(
        R2_SB_SB3_n819), .A4(R2_SB_SB3_n818), .ZN(R2_SB_SB3_n822) );
  INV_X1 R2_SB_SB3_U229 ( .A(R2_SB_SB3_n789), .ZN(R2_SB_SB3_n853) );
  NOR2_X1 R2_SB_SB3_U228 ( .A1(R2_SB_SB3_n743), .A2(R2_SB_SB3_n603), .ZN(
        R2_SB_SB3_n718) );
  AOI221_X1 R2_SB_SB3_U227 ( .B1(R2_SB_SB3_n877), .B2(R2_SB_SB3_n684), .C1(
        R2_SB_SB3_n591), .C2(R2_SB_SB3_n89), .A(R2_SB_SB3_n590), .ZN(
        R2_SB_SB3_n593) );
  AOI22_X1 R2_SB_SB3_U226 ( .A1(R2_SB_SB3_n810), .A2(R2_SB_SB3_n589), .B1(
        R2_SB_SB3_n798), .B2(R2_SB_SB3_n723), .ZN(R2_SB_SB3_n594) );
  OAI221_X1 R2_SB_SB3_U225 ( .B1(R2_SB_SB3_n594), .B2(R2_SB_SB3_n859), .C1(
        R2_SB_SB3_n593), .C2(R2_SB_SB3_n849), .A(R2_SB_SB3_n592), .ZN(
        R2_SB_SB3_n596) );
  INV_X1 R2_SB_SB3_U224 ( .A(R2_SB_SB3_n744), .ZN(R2_SB_SB3_n868) );
  OAI21_X1 R2_SB_SB3_U223 ( .B1(R2_SB_SB3_n779), .B2(R2_SB_SB3_n453), .A(
        R2_SB_SB3_n656), .ZN(R2_SB_SB3_n503) );
  NOR2_X1 R2_SB_SB3_U222 ( .A1(R2_SB_SB3_n618), .A2(R2_SB_SB3_n780), .ZN(
        R2_SB_SB3_n504) );
  OAI221_X1 R2_SB_SB3_U221 ( .B1(R2_SB_SB3_n504), .B2(R2_SB_SB3_n840), .C1(
        R2_SB_SB3_n869), .C2(R2_SB_SB3_n852), .A(R2_SB_SB3_n503), .ZN(
        R2_SB_SB3_n505) );
  INV_X1 R2_SB_SB3_U220 ( .A(R2_SB_SB3_n617), .ZN(R2_SB_SB3_n862) );
  AOI21_X1 R2_SB_SB3_U219 ( .B1(R2_SB_SB3_n828), .B2(R2_SB_SB3_n850), .A(
        R2_SB_SB3_n879), .ZN(R2_SB_SB3_n459) );
  AOI221_X1 R2_SB_SB3_U218 ( .B1(R2_SB_SB3_n463), .B2(R2_SB_SB3_n591), .C1(
        R2_SB_SB3_n514), .C2(R2_SB_SB3_n766), .A(R2_SB_SB3_n459), .ZN(
        R2_SB_SB3_n488) );
  OAI222_X1 R2_SB_SB3_U217 ( .A1(R2_SB_SB3_n623), .A2(R2_SB_SB3_n851), .B1(
        R2_SB_SB3_n622), .B2(R2_SB_SB3_n883), .C1(R2_SB_SB3_n621), .C2(
        R2_SB_SB3_n905), .ZN(R2_SB_SB3_n624) );
  OAI221_X1 R2_SB_SB3_U216 ( .B1(R2_SB_SB3_n903), .B2(R2_SB_SB3_n844), .C1(
        R2_SB_SB3_n848), .C2(R2_SB_SB3_n910), .A(R2_SB_SB3_n607), .ZN(
        R2_SB_SB3_n626) );
  OAI211_X1 R2_SB_SB3_U215 ( .C1(R2_SB_SB3_n857), .C2(R2_SB_SB3_n831), .A(
        R2_SB_SB3_n612), .B(R2_SB_SB3_n611), .ZN(R2_SB_SB3_n625) );
  AOI221_X1 R2_SB_SB3_U214 ( .B1(R2_SB_SB3_n452), .B2(R2_SB_SB3_n626), .C1(
        R2_SB_SB3_n752), .C2(R2_SB_SB3_n625), .A(R2_SB_SB3_n624), .ZN(
        R2_SB_SB3_n644) );
  OAI22_X1 R2_SB_SB3_U213 ( .A1(R2_SB_SB3_n733), .A2(R2_SB_SB3_n837), .B1(
        R2_SB_SB3_n842), .B2(R2_SB_SB3_n884), .ZN(R2_SB_SB3_n653) );
  OAI22_X1 R2_SB_SB3_U212 ( .A1(R2_SB_SB3_n858), .A2(R2_SB_SB3_n834), .B1(
        R2_SB_n306), .B2(R2_SB_SB3_n859), .ZN(R2_SB_SB3_n654) );
  OAI21_X1 R2_SB_SB3_U211 ( .B1(R2_SB_SB3_n903), .B2(R2_SB_SB3_n859), .A(
        R2_SB_SB3_n895), .ZN(R2_SB_SB3_n655) );
  AOI221_X1 R2_SB_SB3_U210 ( .B1(R2_SB_SB3_n795), .B2(R2_SB_SB3_n655), .C1(
        R2_SB_SB3_n702), .C2(R2_SB_SB3_n654), .A(R2_SB_SB3_n653), .ZN(
        R2_SB_SB3_n692) );
  AOI221_X1 R2_SB_SB3_U209 ( .B1(R2_SB_SB3_n684), .B2(R2_SB_SB3_n536), .C1(
        R2_SB_SB3_n535), .C2(R2_SB_SB3_n628), .A(R2_SB_SB3_n534), .ZN(
        R2_SB_SB3_n537) );
  OAI222_X1 R2_SB_SB3_U208 ( .A1(R2_SB_SB3_n543), .A2(R2_SB_SB3_n847), .B1(
        R2_SB_SB3_n835), .B2(R2_SB_SB3_n573), .C1(R2_SB_SB3_n542), .C2(
        R2_SB_SB3_n883), .ZN(R2_SB_SB3_n544) );
  OAI221_X1 R2_SB_SB3_U207 ( .B1(R2_SB_SB3_n89), .B2(R2_SB_SB3_n588), .C1(
        R2_SB_n305), .C2(R2_SB_SB3_n910), .A(R2_SB_SB3_n537), .ZN(
        R2_SB_SB3_n545) );
  AOI221_X1 R2_SB_SB3_U206 ( .B1(R2_SB_SB3_n792), .B2(R2_SB_SB3_n545), .C1(
        R2_SB_SB3_n753), .C2(R2_SB_SB3_n791), .A(R2_SB_SB3_n544), .ZN(
        R2_SB_SB3_n560) );
  AOI22_X1 R2_SB_SB3_U205 ( .A1(R2_SB_SB3_n798), .A2(R2_SB_SB3_n708), .B1(
        R2_SB_SB3_n795), .B2(R2_SB_SB3_n767), .ZN(R2_SB_SB3_n631) );
  AOI21_X1 R2_SB_SB3_U204 ( .B1(R2_SB_SB3_n755), .B2(R2_SB_SB3_n758), .A(
        R2_SB_SB3_n756), .ZN(R2_SB_SB3_n629) );
  OAI222_X1 R2_SB_SB3_U203 ( .A1(R2_SB_SB3_n631), .A2(R2_SB_SB3_n857), .B1(
        R2_SB_SB3_n630), .B2(R2_SB_SB3_n875), .C1(R2_SB_n306), .C2(
        R2_SB_SB3_n629), .ZN(R2_SB_SB3_n632) );
  AOI221_X1 R2_SB_SB3_U202 ( .B1(R2_SB_SB3_n725), .B2(R2_SB_SB3_n728), .C1(
        R2_SB_SB3_n651), .C2(R2_SB_SB3_n789), .A(R2_SB_SB3_n632), .ZN(
        R2_SB_SB3_n643) );
  OAI222_X1 R2_SB_SB3_U201 ( .A1(R2_SB_SB3_n865), .A2(R2_SB_SB3_n785), .B1(
        R2_SB_SB3_n784), .B2(R2_SB_SB3_n905), .C1(R2_SB_SB3_n827), .C2(
        R2_SB_SB3_n897), .ZN(R2_SB_SB3_n786) );
  OAI211_X1 R2_SB_SB3_U200 ( .C1(R2_SB_SB3_n829), .C2(R2_SB_SB3_n770), .A(
        R2_SB_SB3_n769), .B(R2_SB_SB3_n768), .ZN(R2_SB_SB3_n788) );
  OAI211_X1 R2_SB_SB3_U199 ( .C1(R2_SB_SB3_n895), .C2(R2_SB_SB3_n848), .A(
        R2_SB_SB3_n777), .B(R2_SB_SB3_n887), .ZN(R2_SB_SB3_n787) );
  AOI221_X1 R2_SB_SB3_U198 ( .B1(R2_SB_SB3_n789), .B2(R2_SB_SB3_n788), .C1(
        R2_SB_n305), .C2(R2_SB_SB3_n787), .A(R2_SB_SB3_n786), .ZN(
        R2_SB_SB3_n823) );
  INV_X1 R2_SB_SB3_U197 ( .A(R2_SB_SB3_n656), .ZN(R2_SB_SB3_n859) );
  AOI211_X1 R2_SB_SB3_U196 ( .C1(R2_SB_SB3_n789), .C2(R2_SB_SB3_n812), .A(
        R2_SB_SB3_n882), .B(R2_SB_SB3_n727), .ZN(R2_SB_SB3_n577) );
  AOI211_X1 R2_SB_SB3_U195 ( .C1(R2_SB_SB3_n744), .C2(R2_SB_SB3_n843), .A(
        R2_SB_SB3_n730), .B(R2_SB_SB3_n792), .ZN(R2_SB_SB3_n509) );
  AOI21_X1 R2_SB_SB3_U194 ( .B1(R2_SB_SB3_n854), .B2(R2_SB_SB3_n881), .A(
        R2_SB_SB3_n767), .ZN(R2_SB_SB3_n477) );
  OAI222_X1 R2_SB_SB3_U193 ( .A1(R2_SB_SB3_n843), .A2(R2_SB_SB3_n885), .B1(
        R2_SB_SB3_n477), .B2(R2_SB_SB3_n845), .C1(R2_SB_SB3_n864), .C2(
        R2_SB_SB3_n878), .ZN(R2_SB_SB3_n479) );
  OAI22_X1 R2_SB_SB3_U192 ( .A1(R2_SB_SB3_n849), .A2(R2_SB_SB3_n648), .B1(
        R2_SB_SB3_n862), .B2(R2_SB_SB3_n844), .ZN(R2_SB_SB3_n478) );
  AOI211_X1 R2_SB_SB3_U191 ( .C1(R2_SB_SB3_n791), .C2(R2_SB_SB3_n812), .A(
        R2_SB_SB3_n479), .B(R2_SB_SB3_n478), .ZN(R2_SB_SB3_n480) );
  NOR3_X1 R2_SB_SB3_U190 ( .A1(R2_SB_SB3_n838), .A2(R2_SB_n305), .A3(
        R2_SB_SB3_n864), .ZN(R2_SB_SB3_n610) );
  AOI21_X1 R2_SB_SB3_U189 ( .B1(R2_SB_SB3_n858), .B2(R2_SB_SB3_n608), .A(
        R2_SB_SB3_n827), .ZN(R2_SB_SB3_n609) );
  AOI211_X1 R2_SB_SB3_U188 ( .C1(R2_SB_SB3_n646), .C2(R2_SB_SB3_n781), .A(
        R2_SB_SB3_n610), .B(R2_SB_SB3_n609), .ZN(R2_SB_SB3_n611) );
  INV_X1 R2_SB_SB3_U187 ( .A(R2_SB_SB3_n752), .ZN(R2_SB_SB3_n878) );
  NOR2_X1 R2_SB_SB3_U186 ( .A1(R2_SB_SB3_n857), .A2(R2_SB_SB3_n863), .ZN(
        R2_SB_SB3_n670) );
  INV_X1 R2_SB_SB3_U185 ( .A(R2_SB_SB3_n772), .ZN(R2_SB_SB3_n883) );
  INV_X1 R2_SB_SB3_U184 ( .A(R2_SB_SB3_n618), .ZN(R2_SB_SB3_n864) );
  OAI21_X1 R2_SB_SB3_U183 ( .B1(R2_SB_SB3_n856), .B2(R2_SB_SB3_n874), .A(
        R2_SB_SB3_n893), .ZN(R2_SB_SB3_n516) );
  AOI21_X1 R2_SB_SB3_U182 ( .B1(R2_SB_SB3_n781), .B2(R2_SB_SB3_n516), .A(
        R2_SB_SB3_n515), .ZN(R2_SB_SB3_n517) );
  AOI21_X1 R2_SB_SB3_U181 ( .B1(R2_SB_SB3_n900), .B2(R2_SB_SB3_n603), .A(
        R2_SB_SB3_n783), .ZN(R2_SB_SB3_n518) );
  OAI221_X1 R2_SB_SB3_U180 ( .B1(R2_SB_SB3_n518), .B2(R2_SB_SB3_n453), .C1(
        R2_SB_SB3_n838), .C2(R2_SB_SB3_n904), .A(R2_SB_SB3_n517), .ZN(
        R2_SB_SB3_n523) );
  AOI21_X1 R2_SB_SB3_U179 ( .B1(R2_SB_SB3_n646), .B2(R2_SB_SB3_n634), .A(
        R2_SB_SB3_n633), .ZN(R2_SB_SB3_n636) );
  OAI21_X1 R2_SB_SB3_U178 ( .B1(R2_SB_SB3_n747), .B2(R2_SB_SB3_n799), .A(
        R2_SB_SB3_n882), .ZN(R2_SB_SB3_n635) );
  NAND2_X1 R2_SB_SB3_U177 ( .A1(R2_SB_SB3_n828), .A2(R2_SB_SB3_n843), .ZN(
        R2_SB_SB3_n637) );
  OAI221_X1 R2_SB_SB3_U176 ( .B1(R2_SB_SB3_n910), .B2(R2_SB_SB3_n637), .C1(
        R2_SB_SB3_n636), .C2(R2_SB_SB3_n829), .A(R2_SB_SB3_n635), .ZN(
        R2_SB_SB3_n641) );
  OAI22_X1 R2_SB_SB3_U175 ( .A1(R2_SB_SB3_n857), .A2(R2_SB_SB3_n838), .B1(
        R2_SB_SB3_n832), .B2(R2_SB_SB3_n865), .ZN(R2_SB_SB3_n469) );
  OAI21_X1 R2_SB_SB3_U174 ( .B1(R2_SB_n306), .B2(R2_SB_SB3_n845), .A(
        R2_SB_SB3_n849), .ZN(R2_SB_SB3_n471) );
  AOI221_X1 R2_SB_SB3_U173 ( .B1(R2_SB_SB3_n744), .B2(R2_SB_SB3_n471), .C1(
        R2_SB_SB3_n470), .C2(R2_SB_SB3_n863), .A(R2_SB_SB3_n469), .ZN(
        R2_SB_SB3_n476) );
  AOI221_X1 R2_SB_SB3_U172 ( .B1(R2_SB_SB3_n882), .B2(R2_SB_SB3_n792), .C1(
        R2_SB_SB3_n627), .C2(R2_SB_SB3_n702), .A(R2_SB_SB3_n698), .ZN(
        R2_SB_SB3_n583) );
  NOR2_X1 R2_SB_SB3_U171 ( .A1(R2_SB_SB3_n813), .A2(R2_SB_SB3_n694), .ZN(
        R2_SB_SB3_n695) );
  OAI221_X1 R2_SB_SB3_U170 ( .B1(R2_SB_SB3_n695), .B2(R2_SB_SB3_n851), .C1(
        R2_SB_SB3_n856), .C2(R2_SB_SB3_n878), .A(R2_SB_SB3_n904), .ZN(
        R2_SB_SB3_n697) );
  INV_X1 R2_SB_SB3_U169 ( .A(R2_SB_SB3_n801), .ZN(R2_SB_SB3_n873) );
  AOI222_X1 R2_SB_SB3_U168 ( .A1(R2_SB_SB3_n771), .A2(R2_SB_SB3_n698), .B1(
        R2_SB_SB3_n781), .B2(R2_SB_SB3_n697), .C1(R2_SB_SB3_n696), .C2(
        R2_SB_SB3_n873), .ZN(R2_SB_SB3_n741) );
  AOI22_X1 R2_SB_SB3_U167 ( .A1(R2_SB_SB3_n758), .A2(R2_SB_SB3_n694), .B1(
        R2_SB_SB3_n779), .B2(R2_SB_SB3_n863), .ZN(R2_SB_SB3_n619) );
  OAI222_X1 R2_SB_SB3_U166 ( .A1(R2_SB_SB3_n864), .A2(R2_SB_SB3_n833), .B1(
        R2_SB_n305), .B2(R2_SB_SB3_n619), .C1(R2_SB_SB3_n858), .C2(
        R2_SB_SB3_n839), .ZN(R2_SB_SB3_n620) );
  AOI221_X1 R2_SB_SB3_U165 ( .B1(R2_SB_SB3_n789), .B2(R2_SB_SB3_n628), .C1(
        R2_SB_SB3_n778), .C2(R2_SB_SB3_n771), .A(R2_SB_SB3_n620), .ZN(
        R2_SB_SB3_n621) );
  NAND2_X1 R2_SB_SB3_U164 ( .A1(R2_SB_SB3_n848), .A2(R2_SB_SB3_n841), .ZN(
        R2_SB_SB3_n616) );
  INV_X1 R2_SB_SB3_U163 ( .A(R2_SB_SB3_n615), .ZN(R2_SB_SB3_n861) );
  AOI221_X1 R2_SB_SB3_U162 ( .B1(R2_SB_SB3_n747), .B2(R2_SB_SB3_n618), .C1(
        R2_SB_SB3_n617), .C2(R2_SB_SB3_n616), .A(R2_SB_SB3_n861), .ZN(
        R2_SB_SB3_n622) );
  OAI221_X1 R2_SB_SB3_U161 ( .B1(R2_SB_SB3_n870), .B2(R2_SB_SB3_n838), .C1(
        R2_SB_SB3_n840), .C2(R2_SB_SB3_n868), .A(R2_SB_SB3_n496), .ZN(
        R2_SB_SB3_n497) );
  OAI211_X1 R2_SB_SB3_U160 ( .C1(R2_SB_SB3_n879), .C2(R2_SB_SB3_n844), .A(
        R2_SB_SB3_n711), .B(R2_SB_SB3_n491), .ZN(R2_SB_SB3_n499) );
  AOI222_X1 R2_SB_SB3_U159 ( .A1(R2_SB_SB3_n499), .A2(R2_SB_SB3_n453), .B1(
        R2_SB_SB3_n498), .B2(R2_SB_SB3_n854), .C1(R2_SB_SB3_n752), .C2(
        R2_SB_SB3_n497), .ZN(R2_SB_SB3_n527) );
  OAI222_X1 R2_SB_SB3_U158 ( .A1(R2_SB_SB3_n865), .A2(R2_SB_SB3_n838), .B1(
        R2_SB_SB3_n699), .B2(R2_SB_SB3_n868), .C1(R2_SB_n306), .C2(
        R2_SB_SB3_n858), .ZN(R2_SB_SB3_n704) );
  OAI22_X1 R2_SB_SB3_U157 ( .A1(R2_SB_SB3_n864), .A2(R2_SB_SB3_n839), .B1(
        R2_SB_SB3_n700), .B2(R2_SB_SB3_n833), .ZN(R2_SB_SB3_n701) );
  AOI222_X1 R2_SB_SB3_U156 ( .A1(R2_SB_SB3_n772), .A2(R2_SB_SB3_n704), .B1(
        R2_SB_SB3_n882), .B2(R2_SB_SB3_n703), .C1(R2_SB_SB3_n702), .C2(
        R2_SB_SB3_n701), .ZN(R2_SB_SB3_n740) );
  NOR2_X1 R2_SB_SB3_U155 ( .A1(R2_SB_SB3_n881), .A2(R2_SB_SB3_n863), .ZN(
        R2_SB_SB3_n634) );
  OAI222_X1 R2_SB_SB3_U154 ( .A1(R2_SB_n306), .A2(R2_SB_SB3_n875), .B1(
        R2_SB_SB3_n883), .B2(R2_SB_SB3_n826), .C1(R2_SB_SB3_n905), .C2(
        R2_SB_SB3_n831), .ZN(R2_SB_SB3_n707) );
  AOI211_X1 R2_SB_SB3_U153 ( .C1(R2_SB_SB3_n709), .C2(R2_SB_SB3_n708), .A(
        R2_SB_SB3_n707), .B(R2_SB_SB3_n706), .ZN(R2_SB_SB3_n710) );
  OAI222_X1 R2_SB_SB3_U152 ( .A1(R2_SB_SB3_n833), .A2(R2_SB_SB3_n898), .B1(
        R2_SB_SB3_n710), .B2(R2_SB_SB3_n859), .C1(R2_SB_SB3_n832), .C2(
        R2_SB_SB3_n800), .ZN(R2_SB_SB3_n712) );
  INV_X1 R2_SB_SB3_U151 ( .A(R2_SB_SB3_n792), .ZN(R2_SB_SB3_n845) );
  OAI221_X1 R2_SB_SB3_U150 ( .B1(R2_SB_SB3_n833), .B2(R2_SB_SB3_n774), .C1(
        R2_SB_SB3_n509), .C2(R2_SB_SB3_n829), .A(R2_SB_SB3_n508), .ZN(
        R2_SB_SB3_n510) );
  AOI221_X1 R2_SB_SB3_U149 ( .B1(R2_SB_SB3_n507), .B2(R2_SB_SB3_n506), .C1(
        R2_SB_SB3_n780), .C2(R2_SB_SB3_n684), .A(R2_SB_SB3_n505), .ZN(
        R2_SB_SB3_n512) );
  AOI221_X1 R2_SB_SB3_U148 ( .B1(R2_SB_SB3_n743), .B2(R2_SB_SB3_n684), .C1(
        R2_SB_SB3_n780), .C2(R2_SB_SB3_n627), .A(R2_SB_SB3_n510), .ZN(
        R2_SB_SB3_n511) );
  OAI222_X1 R2_SB_SB3_U147 ( .A1(R2_SB_SB3_n512), .A2(R2_SB_SB3_n905), .B1(
        R2_SB_SB3_n511), .B2(R2_SB_SB3_n883), .C1(R2_SB_SB3_n884), .C2(
        R2_SB_SB3_n844), .ZN(R2_SB_SB3_n513) );
  INV_X1 R2_SB_SB3_U146 ( .A(R2_SB_SB3_n659), .ZN(R2_SB_SB3_n867) );
  AOI221_X1 R2_SB_SB3_U145 ( .B1(R2_SB_SB3_n794), .B2(R2_SB_SB3_n730), .C1(
        R2_SB_SB3_n742), .C2(R2_SB_SB3_n780), .A(R2_SB_SB3_n867), .ZN(
        R2_SB_SB3_n574) );
  NOR4_X1 R2_SB_SB3_U144 ( .A1(R2_SB_SB3_n452), .A2(R2_SB_SB3_n872), .A3(
        R2_SB_SB3_n849), .A4(R2_SB_SB3_n862), .ZN(R2_SB_SB3_n640) );
  NOR2_X1 R2_SB_SB3_U143 ( .A1(R2_SB_SB3_n89), .A2(R2_SB_SB3_n843), .ZN(
        R2_SB_SB3_n603) );
  NOR2_X1 R2_SB_SB3_U142 ( .A1(R2_SB_SB3_n872), .A2(R2_SB_SB3_n863), .ZN(
        R2_SB_SB3_n812) );
  NOR2_X1 R2_SB_SB3_U141 ( .A1(R2_SB_SB3_n863), .A2(R2_SB_SB3_n854), .ZN(
        R2_SB_SB3_n507) );
  AOI222_X1 R2_SB_SB3_U140 ( .A1(R2_SB_SB3_n782), .A2(R2_SB_SB3_n781), .B1(
        R2_SB_SB3_n780), .B2(R2_SB_SB3_n779), .C1(R2_SB_SB3_n778), .C2(
        R2_SB_SB3_n791), .ZN(R2_SB_SB3_n784) );
  INV_X1 R2_SB_SB3_U139 ( .A(R2_SB_SB3_n795), .ZN(R2_SB_SB3_n838) );
  AOI22_X1 R2_SB_SB3_U138 ( .A1(R2_SB_SB3_n724), .A2(R2_SB_SB3_n810), .B1(
        R2_SB_SB3_n744), .B2(R2_SB_SB3_n723), .ZN(R2_SB_SB3_n726) );
  INV_X1 R2_SB_SB3_U137 ( .A(R2_SB_SB3_n722), .ZN(R2_SB_SB3_n896) );
  INV_X1 R2_SB_SB3_U136 ( .A(R2_SB_SB3_n725), .ZN(R2_SB_SB3_n846) );
  OAI222_X1 R2_SB_SB3_U135 ( .A1(R2_SB_SB3_n849), .A2(R2_SB_SB3_n896), .B1(
        R2_SB_SB3_n726), .B2(R2_SB_SB3_n878), .C1(R2_SB_SB3_n846), .C2(
        R2_SB_SB3_n910), .ZN(R2_SB_SB3_n735) );
  OAI222_X1 R2_SB_SB3_U134 ( .A1(R2_SB_SB3_n853), .A2(R2_SB_SB3_n829), .B1(
        R2_SB_SB3_n608), .B2(R2_SB_SB3_n826), .C1(R2_SB_SB3_n870), .C2(
        R2_SB_SB3_n831), .ZN(R2_SB_SB3_n465) );
  NOR3_X1 R2_SB_SB3_U133 ( .A1(R2_SB_SB3_n877), .A2(R2_SB_SB3_n638), .A3(
        R2_SB_SB3_n679), .ZN(R2_SB_SB3_n466) );
  INV_X1 R2_SB_SB3_U132 ( .A(R2_SB_SB3_n465), .ZN(R2_SB_SB3_n871) );
  OAI222_X1 R2_SB_SB3_U131 ( .A1(R2_SB_SB3_n871), .A2(R2_SB_SB3_n883), .B1(
        R2_SB_SB3_n849), .B2(R2_SB_SB3_n769), .C1(R2_SB_SB3_n466), .C2(
        R2_SB_SB3_n834), .ZN(R2_SB_SB3_n484) );
  INV_X1 R2_SB_SB3_U130 ( .A(R2_SB_SB3_n782), .ZN(R2_SB_SB3_n849) );
  NOR2_X1 R2_SB_SB3_U129 ( .A1(R2_SB_SB3_n830), .A2(R2_SB_SB3_n854), .ZN(
        R2_SB_SB3_n627) );
  NOR2_X1 R2_SB_SB3_U128 ( .A1(R2_SB_SB3_n881), .A2(R2_SB_SB3_n872), .ZN(
        R2_SB_SB3_n669) );
  INV_X1 R2_SB_SB3_U127 ( .A(R2_SB_SB3_n702), .ZN(R2_SB_SB3_n905) );
  NOR2_X1 R2_SB_SB3_U126 ( .A1(R2_SB_SB3_n453), .A2(R2_SB_SB3_n830), .ZN(
        R2_SB_SB3_n766) );
  NOR3_X1 R2_SB_SB3_U125 ( .A1(R2_SB_SB3_n828), .A2(R2_SB_SB3_n854), .A3(
        R2_SB_SB3_n908), .ZN(R2_SB_SB3_n673) );
  NOR2_X1 R2_SB_SB3_U124 ( .A1(R2_SB_SB3_n89), .A2(R2_SB_SB3_n830), .ZN(
        R2_SB_SB3_n771) );
  NOR2_X1 R2_SB_SB3_U123 ( .A1(R2_SB_SB3_n863), .A2(R2_SB_SB3_n843), .ZN(
        R2_SB_SB3_n778) );
  NOR2_X1 R2_SB_SB3_U122 ( .A1(R2_SB_SB3_n830), .A2(R2_SB_n306), .ZN(
        R2_SB_SB3_n779) );
  AOI21_X1 R2_SB_SB3_U121 ( .B1(R2_SB_SB3_n826), .B2(R2_SB_SB3_n833), .A(
        R2_SB_SB3_n800), .ZN(R2_SB_SB3_n549) );
  INV_X1 R2_SB_SB3_U120 ( .A(R2_SB_SB3_n549), .ZN(R2_SB_SB3_n902) );
  AND3_X1 R2_SB_SB3_U119 ( .A1(R2_SB_SB3_n548), .A2(R2_SB_SB3_n838), .A3(
        R2_SB_SB3_n849), .ZN(R2_SB_SB3_n550) );
  OR3_X1 R2_SB_SB3_U118 ( .A1(R2_SB_SB3_n864), .A2(R2_SB_SB3_n814), .A3(
        R2_SB_SB3_n890), .ZN(R2_SB_SB3_n815) );
  INV_X1 R2_SB_SB3_U117 ( .A(R2_SB_SB3_n519), .ZN(R2_SB_SB3_n886) );
  INV_X1 R2_SB_SB3_U116 ( .A(R2_SB_SB3_n790), .ZN(R2_SB_SB3_n866) );
  NAND2_X1 R2_SB_SB3_U115 ( .A1(R2_SB_SB3_n874), .A2(R2_SB_SB3_n901), .ZN(
        R2_SB_SB3_n728) );
  NAND2_X1 R2_SB_SB3_U114 ( .A1(R2_SB_SB3_n890), .A2(R2_SB_SB3_n874), .ZN(
        R2_SB_SB3_n536) );
  NAND2_X1 R2_SB_SB3_U113 ( .A1(R2_SB_SB3_n836), .A2(R2_SB_SB3_n826), .ZN(
        R2_SB_SB3_n723) );
  NAND2_X1 R2_SB_SB3_U112 ( .A1(R2_SB_SB3_n905), .A2(R2_SB_SB3_n875), .ZN(
        R2_SB_SB3_n589) );
  INV_X1 R2_SB_SB3_U111 ( .A(R2_SB_SB3_n627), .ZN(R2_SB_SB3_n856) );
  NAND2_X1 R2_SB_SB3_U110 ( .A1(R2_SB_SB3_n836), .A2(R2_SB_SB3_n829), .ZN(
        R2_SB_SB3_n748) );
  AND2_X1 R2_SB_SB3_U109 ( .A1(R2_SB_SB3_n766), .A2(R2_SB_SB3_n671), .ZN(
        R2_SB_SB3_n555) );
  INV_X1 R2_SB_SB3_U108 ( .A(R2_SB_SB3_n812), .ZN(R2_SB_SB3_n875) );
  OAI21_X1 R2_SB_SB3_U107 ( .B1(R2_SB_SB3_n847), .B2(R2_SB_SB3_n895), .A(
        R2_SB_SB3_n800), .ZN(R2_SB_SB3_n806) );
  NAND2_X1 R2_SB_SB3_U106 ( .A1(R2_SB_SB3_n628), .A2(R2_SB_SB3_n634), .ZN(
        R2_SB_SB3_n769) );
  NAND2_X1 R2_SB_SB3_U105 ( .A1(R2_SB_SB3_n507), .A2(R2_SB_SB3_n669), .ZN(
        R2_SB_SB3_n588) );
  INV_X1 R2_SB_SB3_U104 ( .A(R2_SB_SB3_n634), .ZN(R2_SB_SB3_n903) );
  INV_X1 R2_SB_SB3_U103 ( .A(R2_SB_SB3_n778), .ZN(R2_SB_SB3_n865) );
  NOR2_X1 R2_SB_SB3_U102 ( .A1(R2_SB_SB3_n730), .A2(R2_SB_SB3_n758), .ZN(
        R2_SB_SB3_n685) );
  AOI21_X1 R2_SB_SB3_U101 ( .B1(R2_SB_SB3_n588), .B2(R2_SB_SB3_n773), .A(
        R2_SB_SB3_n836), .ZN(R2_SB_SB3_n460) );
  AOI21_X1 R2_SB_SB3_U100 ( .B1(R2_SB_SB3_n802), .B2(R2_SB_SB3_n801), .A(
        R2_SB_SB3_n835), .ZN(R2_SB_SB3_n803) );
  INV_X1 R2_SB_SB3_U99 ( .A(R2_SB_SB3_n672), .ZN(R2_SB_SB3_n888) );
  NOR4_X1 R2_SB_SB3_U98 ( .A1(R2_SB_SB3_n675), .A2(R2_SB_SB3_n888), .A3(
        R2_SB_SB3_n674), .A4(R2_SB_SB3_n673), .ZN(R2_SB_SB3_n676) );
  NAND2_X1 R2_SB_SB3_U97 ( .A1(R2_SB_SB3_n778), .A2(R2_SB_SB3_n669), .ZN(
        R2_SB_SB3_n573) );
  INV_X1 R2_SB_SB3_U96 ( .A(R2_SB_SB3_n648), .ZN(R2_SB_SB3_n882) );
  NOR2_X1 R2_SB_SB3_U95 ( .A1(R2_SB_SB3_n849), .A2(R2_SB_SB3_n89), .ZN(
        R2_SB_SB3_n502) );
  NOR2_X1 R2_SB_SB3_U94 ( .A1(R2_SB_SB3_n851), .A2(R2_SB_n306), .ZN(
        R2_SB_SB3_n470) );
  NOR2_X1 R2_SB_SB3_U93 ( .A1(R2_SB_SB3_n853), .A2(R2_SB_SB3_n903), .ZN(
        R2_SB_SB3_n514) );
  INV_X1 R2_SB_SB3_U92 ( .A(R2_SB_SB3_n604), .ZN(R2_SB_SB3_n844) );
  NOR2_X1 R2_SB_SB3_U91 ( .A1(R2_SB_SB3_n862), .A2(R2_SB_SB3_n883), .ZN(
        R2_SB_SB3_n534) );
  INV_X1 R2_SB_SB3_U90 ( .A(R2_SB_SB3_n603), .ZN(R2_SB_SB3_n848) );
  INV_X1 R2_SB_SB3_U89 ( .A(R2_SB_SB3_n802), .ZN(R2_SB_SB3_n877) );
  NOR2_X1 R2_SB_SB3_U88 ( .A1(R2_SB_SB3_n905), .A2(R2_SB_SB3_n866), .ZN(
        R2_SB_SB3_n671) );
  OAI22_X1 R2_SB_SB3_U87 ( .A1(R2_SB_SB3_n730), .A2(R2_SB_SB3_n905), .B1(
        R2_SB_SB3_n901), .B2(R2_SB_SB3_n851), .ZN(R2_SB_SB3_n462) );
  OAI22_X1 R2_SB_SB3_U86 ( .A1(R2_SB_SB3_n875), .A2(R2_SB_SB3_n833), .B1(
        R2_SB_SB3_n874), .B2(R2_SB_SB3_n832), .ZN(R2_SB_SB3_n804) );
  OAI22_X1 R2_SB_SB3_U85 ( .A1(R2_SB_SB3_n665), .A2(R2_SB_SB3_n892), .B1(
        R2_SB_SB3_n841), .B2(R2_SB_SB3_n801), .ZN(R2_SB_SB3_n666) );
  INV_X1 R2_SB_SB3_U84 ( .A(R2_SB_SB3_n758), .ZN(R2_SB_SB3_n847) );
  AOI21_X1 R2_SB_SB3_U83 ( .B1(R2_SB_SB3_n868), .B2(R2_SB_SB3_n845), .A(
        R2_SB_SB3_n785), .ZN(R2_SB_SB3_n687) );
  OAI22_X1 R2_SB_SB3_U82 ( .A1(R2_SB_SB3_n831), .A2(R2_SB_SB3_n895), .B1(
        R2_SB_n305), .B2(R2_SB_SB3_n648), .ZN(R2_SB_SB3_n532) );
  AOI22_X1 R2_SB_SB3_U81 ( .A1(R2_SB_SB3_n758), .A2(R2_SB_n306), .B1(
        R2_SB_SB3_n771), .B2(R2_SB_SB3_n452), .ZN(R2_SB_SB3_n699) );
  INV_X1 R2_SB_SB3_U80 ( .A(R2_SB_SB3_n771), .ZN(R2_SB_SB3_n831) );
  NOR2_X1 R2_SB_SB3_U79 ( .A1(R2_SB_SB3_n842), .A2(R2_SB_SB3_n898), .ZN(
        R2_SB_SB3_n675) );
  NOR2_X1 R2_SB_SB3_U78 ( .A1(R2_SB_SB3_n868), .A2(R2_SB_SB3_n890), .ZN(
        R2_SB_SB3_n576) );
  NOR2_X1 R2_SB_SB3_U77 ( .A1(R2_SB_SB3_n774), .A2(R2_SB_SB3_n890), .ZN(
        R2_SB_SB3_n565) );
  NOR2_X1 R2_SB_SB3_U76 ( .A1(R2_SB_SB3_n845), .A2(R2_SB_SB3_n89), .ZN(
        R2_SB_SB3_n725) );
  NOR2_X1 R2_SB_SB3_U75 ( .A1(R2_SB_SB3_n853), .A2(R2_SB_SB3_n890), .ZN(
        R2_SB_SB3_n633) );
  NOR2_X1 R2_SB_SB3_U74 ( .A1(R2_SB_SB3_n868), .A2(R2_SB_SB3_n905), .ZN(
        R2_SB_SB3_n754) );
  NOR2_X1 R2_SB_SB3_U73 ( .A1(R2_SB_SB3_n869), .A2(R2_SB_SB3_n905), .ZN(
        R2_SB_SB3_n698) );
  NOR2_X1 R2_SB_SB3_U72 ( .A1(R2_SB_SB3_n898), .A2(R2_SB_SB3_n845), .ZN(
        R2_SB_SB3_n756) );
  NOR2_X1 R2_SB_SB3_U71 ( .A1(R2_SB_SB3_n774), .A2(R2_SB_SB3_n905), .ZN(
        R2_SB_SB3_n638) );
  NOR2_X1 R2_SB_SB3_U70 ( .A1(R2_SB_SB3_n870), .A2(R2_SB_SB3_n890), .ZN(
        R2_SB_SB3_n727) );
  OAI22_X1 R2_SB_SB3_U69 ( .A1(R2_SB_SB3_n453), .A2(R2_SB_SB3_n879), .B1(
        R2_SB_SB3_n89), .B2(R2_SB_SB3_n880), .ZN(R2_SB_SB3_n538) );
  AOI211_X1 R2_SB_SB3_U68 ( .C1(R2_SB_SB3_n576), .C2(R2_SB_SB3_n89), .A(
        R2_SB_SB3_n538), .B(R2_SB_SB3_n722), .ZN(R2_SB_SB3_n543) );
  INV_X1 R2_SB_SB3_U67 ( .A(R2_SB_SB3_n779), .ZN(R2_SB_SB3_n833) );
  NOR3_X1 R2_SB_SB3_U66 ( .A1(R2_SB_SB3_n841), .A2(R2_SB_SB3_n858), .A3(
        R2_SB_SB3_n874), .ZN(R2_SB_SB3_n521) );
  INV_X1 R2_SB_SB3_U65 ( .A(R2_SB_SB3_n766), .ZN(R2_SB_SB3_n835) );
  NOR2_X1 R2_SB_SB3_U64 ( .A1(R2_SB_SB3_n838), .A2(R2_SB_SB3_n453), .ZN(
        R2_SB_SB3_n742) );
  INV_X1 R2_SB_SB3_U63 ( .A(R2_SB_SB3_n730), .ZN(R2_SB_SB3_n858) );
  NOR2_X1 R2_SB_SB3_U62 ( .A1(R2_SB_SB3_n878), .A2(R2_SB_SB3_n869), .ZN(
        R2_SB_SB3_n713) );
  NOR2_X1 R2_SB_SB3_U61 ( .A1(R2_SB_SB3_n833), .A2(R2_SB_SB3_n453), .ZN(
        R2_SB_SB3_n799) );
  AOI22_X1 R2_SB_SB3_U60 ( .A1(R2_SB_SB3_n877), .A2(R2_SB_SB3_n452), .B1(
        R2_SB_SB3_n781), .B2(R2_SB_SB3_n669), .ZN(R2_SB_SB3_n500) );
  OAI211_X1 R2_SB_SB3_U59 ( .C1(R2_SB_SB3_n89), .C2(R2_SB_SB3_n893), .A(
        R2_SB_SB3_n907), .B(R2_SB_SB3_n500), .ZN(R2_SB_SB3_n501) );
  AOI222_X1 R2_SB_SB3_U58 ( .A1(R2_SB_SB3_n591), .A2(R2_SB_SB3_n748), .B1(
        R2_SB_SB3_n502), .B2(R2_SB_SB3_n679), .C1(R2_SB_SB3_n758), .C2(
        R2_SB_SB3_n501), .ZN(R2_SB_SB3_n526) );
  OAI222_X1 R2_SB_SB3_U57 ( .A1(R2_SB_SB3_n845), .A2(R2_SB_SB3_n880), .B1(
        R2_SB_SB3_n835), .B2(R2_SB_SB3_n898), .C1(R2_SB_SB3_n836), .C2(
        R2_SB_SB3_n894), .ZN(R2_SB_SB3_n602) );
  NOR2_X1 R2_SB_SB3_U56 ( .A1(R2_SB_SB3_n883), .A2(R2_SB_SB3_n869), .ZN(
        R2_SB_SB3_n755) );
  NOR2_X1 R2_SB_SB3_U55 ( .A1(R2_SB_SB3_n862), .A2(R2_SB_SB3_n890), .ZN(
        R2_SB_SB3_n753) );
  NOR2_X1 R2_SB_SB3_U54 ( .A1(R2_SB_SB3_n862), .A2(R2_SB_SB3_n905), .ZN(
        R2_SB_SB3_n759) );
  NOR2_X1 R2_SB_SB3_U53 ( .A1(R2_SB_SB3_n862), .A2(R2_SB_SB3_n878), .ZN(
        R2_SB_SB3_n591) );
  NOR2_X1 R2_SB_SB3_U52 ( .A1(R2_SB_SB3_n869), .A2(R2_SB_SB3_n890), .ZN(
        R2_SB_SB3_n679) );
  INV_X1 R2_SB_SB3_U51 ( .A(R2_SB_SB3_n669), .ZN(R2_SB_SB3_n890) );
  NOR2_X2 R2_SB_SB3_U50 ( .A1(R2_SB_SB3_n89), .A2(R2_SB_SB3_n453), .ZN(
        R2_SB_SB3_n781) );
  NOR2_X2 R2_SB_SB3_U49 ( .A1(R2_SB_SB3_n89), .A2(R2_SB_SB3_n452), .ZN(
        R2_SB_SB3_n684) );
  NOR3_X1 R2_SB_SB3_U48 ( .A1(R2_SB_SB3_n878), .A2(R2_SB_SB3_n866), .A3(
        R2_SB_SB3_n838), .ZN(R2_SB_SB3_n674) );
  NOR2_X1 R2_SB_SB3_U47 ( .A1(R2_SB_SB3_n840), .A2(R2_SB_SB3_n452), .ZN(
        R2_SB_SB3_n747) );
  NOR2_X1 R2_SB_SB3_U46 ( .A1(R2_SB_SB3_n453), .A2(R2_SB_n306), .ZN(
        R2_SB_SB3_n810) );
  INV_X1 R2_SB_SB3_U45 ( .A(R2_SB_SB3_n633), .ZN(R2_SB_SB3_n891) );
  INV_X1 R2_SB_SB3_U44 ( .A(R2_SB_SB3_n534), .ZN(R2_SB_SB3_n885) );
  INV_X1 R2_SB_SB3_U43 ( .A(R2_SB_SB3_n470), .ZN(R2_SB_SB3_n852) );
  INV_X1 R2_SB_SB3_U42 ( .A(R2_SB_SB3_n502), .ZN(R2_SB_SB3_n850) );
  INV_X1 R2_SB_SB3_U41 ( .A(R2_SB_SB3_n514), .ZN(R2_SB_SB3_n904) );
  INV_X1 R2_SB_SB3_U40 ( .A(R2_SB_SB3_n698), .ZN(R2_SB_SB3_n906) );
  INV_X1 R2_SB_SB3_U39 ( .A(R2_SB_SB3_n638), .ZN(R2_SB_SB3_n908) );
  INV_X1 R2_SB_SB3_U38 ( .A(R2_SB_SB3_n565), .ZN(R2_SB_SB3_n892) );
  INV_X1 R2_SB_SB3_U37 ( .A(R2_SB_SB3_n753), .ZN(R2_SB_SB3_n893) );
  INV_X1 R2_SB_SB3_U36 ( .A(R2_SB_SB3_n727), .ZN(R2_SB_SB3_n894) );
  INV_X1 R2_SB_SB3_U35 ( .A(R2_SB_SB3_n755), .ZN(R2_SB_SB3_n884) );
  INV_X1 R2_SB_SB3_U34 ( .A(R2_SB_SB3_n799), .ZN(R2_SB_SB3_n834) );
  NAND2_X1 R2_SB_SB3_U33 ( .A1(R2_SB_SB3_n781), .A2(R2_SB_SB3_n671), .ZN(
        R2_SB_SB3_n716) );
  INV_X1 R2_SB_SB3_U32 ( .A(R2_SB_SB3_n588), .ZN(R2_SB_SB3_n900) );
  INV_X1 R2_SB_SB3_U31 ( .A(R2_SB_SB3_n759), .ZN(R2_SB_SB3_n907) );
  INV_X1 R2_SB_SB3_U30 ( .A(R2_SB_SB3_n747), .ZN(R2_SB_SB3_n841) );
  INV_X1 R2_SB_SB3_U29 ( .A(R2_SB_SB3_n713), .ZN(R2_SB_SB3_n879) );
  INV_X1 R2_SB_SB3_U28 ( .A(R2_SB_SB3_n591), .ZN(R2_SB_SB3_n880) );
  INV_X1 R2_SB_SB3_U27 ( .A(R2_SB_SB3_n742), .ZN(R2_SB_SB3_n839) );
  AOI21_X1 R2_SB_SB3_U26 ( .B1(R2_SB_SB3_n848), .B2(R2_SB_SB3_n852), .A(
        R2_SB_SB3_n910), .ZN(R2_SB_SB3_n461) );
  AOI21_X1 R2_SB_SB3_U25 ( .B1(R2_SB_SB3_n831), .B2(R2_SB_SB3_n835), .A(
        R2_SB_SB3_n890), .ZN(R2_SB_SB3_n796) );
  INV_X1 R2_SB_SB3_U24 ( .A(R2_SB_SB3_n684), .ZN(R2_SB_SB3_n827) );
  AOI22_X1 R2_SB_SB3_U23 ( .A1(R2_SB_SB3_n877), .A2(R2_SB_n306), .B1(
        R2_SB_SB3_n713), .B2(R2_SB_SB3_n828), .ZN(R2_SB_SB3_n649) );
  INV_X1 R2_SB_SB3_U22 ( .A(R2_SB_SB3_n754), .ZN(R2_SB_SB3_n910) );
  INV_X1 R2_SB_SB3_U21 ( .A(R2_SB_SB3_n781), .ZN(R2_SB_SB3_n828) );
  INV_X1 R2_SB_SB3_U20 ( .A(R2_SB_SB3_n576), .ZN(R2_SB_SB3_n898) );
  INV_X1 R2_SB_SB3_U19 ( .A(R2_SB_SB3_n679), .ZN(R2_SB_SB3_n895) );
  NOR2_X1 R2_SB_SB3_U18 ( .A1(R2_SB_SB3_n831), .A2(R2_SB_SB3_n452), .ZN(
        R2_SB_SB3_n708) );
  OAI221_X1 R2_SB_SB3_U17 ( .B1(R2_SB_n306), .B2(R2_SB_SB3_n906), .C1(
        R2_SB_SB3_n890), .C2(R2_SB_SB3_n826), .A(R2_SB_SB3_n769), .ZN(
        R2_SB_SB3_n590) );
  NOR2_X1 R2_SB_SB3_U16 ( .A1(R2_SB_SB3_n895), .A2(R2_SB_SB3_n452), .ZN(
        R2_SB_SB3_n722) );
  INV_X1 R2_SB_SB3_U15 ( .A(R2_SB_SB3_n810), .ZN(R2_SB_SB3_n829) );
  NOR2_X1 R2_SB_SB3_U14 ( .A1(R2_SB_n305), .A2(R2_SB_n306), .ZN(R2_SB_SB3_n628) );
  INV_X1 R2_SB_SB3_U13 ( .A(R2_SB_SB3_n708), .ZN(R2_SB_SB3_n832) );
  INV_X1 R2_SB_SB3_U12 ( .A(R2_SB_SB3_n628), .ZN(R2_SB_SB3_n826) );
  NOR2_X1 R2_SB_SB3_U11 ( .A1(R2_SB_SB3_n863), .A2(R2_SB_n309), .ZN(
        R2_SB_SB3_n744) );
  NOR2_X1 R2_SB_SB3_U10 ( .A1(R2_SB_SB3_n881), .A2(R2_SB_n311), .ZN(
        R2_SB_SB3_n772) );
  NOR2_X1 R2_SB_SB3_U9 ( .A1(R2_SB_SB3_n89), .A2(R2_SB_n307), .ZN(
        R2_SB_SB3_n791) );
  NOR2_X1 R2_SB_SB3_U8 ( .A1(R2_SB_SB3_n872), .A2(R2_SB_n312), .ZN(
        R2_SB_SB3_n752) );
  NOR2_X1 R2_SB_SB3_U7 ( .A1(R2_SB_SB3_n854), .A2(R2_SB_SB3_n843), .ZN(
        R2_SB_SB3_n730) );
  NOR2_X1 R2_SB_SB3_U6 ( .A1(R2_SB_SB3_n843), .A2(R2_SB_n310), .ZN(
        R2_SB_SB3_n780) );
  NOR2_X1 R2_SB_SB3_U5 ( .A1(R2_SB_n307), .A2(R2_SB_n308), .ZN(R2_SB_SB3_n743)
         );
  INV_X1 R2_SB_SB3_U4 ( .A(R2_SB_n308), .ZN(R2_SB_SB3_n843) );
  NOR2_X1 R2_SB_SB3_U3 ( .A1(R2_SB_SB3_n453), .A2(R2_SB_n307), .ZN(
        R2_SB_SB3_n696) );
  NOR2_X1 R2_SB_SB3_U2 ( .A1(R2_SB_SB3_n881), .A2(R2_SB_n310), .ZN(
        R2_SB_SB3_n798) );
  NOR2_X1 R2_SB_SB3_U1 ( .A1(R2_SB_SB3_n843), .A2(R2_SB_n309), .ZN(
        R2_SB_SB3_n789) );
  NAND3_X1 R2_SB_SB3_U464 ( .A1(R2_SB_SB3_n772), .A2(R2_SB_SB3_n670), .A3(
        R2_SB_SB3_n794), .ZN(R2_SB_SB3_n519) );
  OAI33_X1 R2_SB_SB3_U463 ( .A1(R2_SB_SB3_n838), .A2(R2_SB_SB3_n858), .A3(
        R2_SB_SB3_n905), .B1(R2_SB_SB3_n853), .B2(R2_SB_SB3_n830), .B3(
        R2_SB_SB3_n874), .ZN(R2_SB_SB3_n467) );
  NAND3_X1 R2_SB_SB3_U462 ( .A1(R2_SB_SB3_n507), .A2(R2_SB_SB3_n702), .A3(
        R2_SB_SB3_n758), .ZN(R2_SB_SB3_n677) );
  OAI33_X1 R2_SB_SB3_U461 ( .A1(R2_SB_SB3_n828), .A2(R2_SB_n312), .A3(
        R2_SB_n307), .B1(R2_SB_SB3_n472), .B2(R2_SB_SB3_n854), .B3(
        R2_SB_SB3_n829), .ZN(R2_SB_SB3_n473) );
  NAND4_X1 R2_SB_SB3_U460 ( .A1(R2_SB_SB3_n488), .A2(R2_SB_SB3_n487), .A3(
        R2_SB_SB3_n486), .A4(R2_SB_SB3_n485), .ZN(R2_SB_n297) );
  NAND3_X1 R2_SB_SB3_U459 ( .A1(R2_SB_SB3_n781), .A2(R2_SB_n307), .A3(
        R2_SB_SB3_n798), .ZN(R2_SB_SB3_n494) );
  NAND4_X1 R2_SB_SB3_U458 ( .A1(R2_SB_SB3_n743), .A2(R2_SB_SB3_n628), .A3(
        R2_SB_SB3_n767), .A4(R2_SB_n312), .ZN(R2_SB_SB3_n493) );
  NAND3_X1 R2_SB_SB3_U457 ( .A1(R2_SB_SB3_n813), .A2(R2_SB_SB3_n830), .A3(
        R2_SB_SB3_n684), .ZN(R2_SB_SB3_n492) );
  NAND3_X1 R2_SB_SB3_U456 ( .A1(R2_SB_SB3_n494), .A2(R2_SB_SB3_n493), .A3(
        R2_SB_SB3_n492), .ZN(R2_SB_SB3_n498) );
  NAND3_X1 R2_SB_SB3_U455 ( .A1(R2_SB_SB3_n844), .A2(R2_SB_SB3_n836), .A3(
        R2_SB_SB3_n548), .ZN(R2_SB_SB3_n506) );
  OAI33_X1 R2_SB_SB3_U454 ( .A1(R2_SB_SB3_n827), .A2(R2_SB_SB3_n856), .A3(
        R2_SB_SB3_n903), .B1(R2_SB_SB3_n898), .B2(R2_SB_SB3_n843), .B3(
        R2_SB_SB3_n826), .ZN(R2_SB_SB3_n515) );
  NAND3_X1 R2_SB_SB3_U453 ( .A1(R2_SB_SB3_n671), .A2(R2_SB_SB3_n453), .A3(
        R2_SB_n307), .ZN(R2_SB_SB3_n816) );
  NAND3_X1 R2_SB_SB3_U452 ( .A1(R2_SB_SB3_n670), .A2(R2_SB_SB3_n669), .A3(
        R2_SB_SB3_n779), .ZN(R2_SB_SB3_n672) );
  NAND3_X1 R2_SB_SB3_U451 ( .A1(R2_SB_SB3_n816), .A2(R2_SB_SB3_n519), .A3(
        R2_SB_SB3_n672), .ZN(R2_SB_SB3_n522) );
  OAI33_X1 R2_SB_SB3_U450 ( .A1(R2_SB_SB3_n832), .A2(R2_SB_SB3_n864), .A3(
        R2_SB_SB3_n890), .B1(R2_SB_SB3_n829), .B2(R2_SB_n312), .B3(
        R2_SB_SB3_n866), .ZN(R2_SB_SB3_n520) );
  NAND4_X1 R2_SB_SB3_U449 ( .A1(R2_SB_SB3_n527), .A2(R2_SB_SB3_n526), .A3(
        R2_SB_SB3_n525), .A4(R2_SB_SB3_n524), .ZN(R2_SB_n298) );
  NAND3_X1 R2_SB_SB3_U448 ( .A1(R2_SB_SB3_n744), .A2(R2_SB_SB3_n603), .A3(
        R2_SB_SB3_n696), .ZN(R2_SB_SB3_n546) );
  NAND3_X1 R2_SB_SB3_U447 ( .A1(R2_SB_SB3_n684), .A2(R2_SB_SB3_n854), .A3(
        R2_SB_SB3_n709), .ZN(R2_SB_SB3_n582) );
  OAI33_X1 R2_SB_SB3_U446 ( .A1(R2_SB_SB3_n859), .A2(R2_SB_SB3_n830), .A3(
        R2_SB_SB3_n901), .B1(R2_SB_SB3_n876), .B2(R2_SB_n306), .B3(
        R2_SB_SB3_n685), .ZN(R2_SB_SB3_n557) );
  NAND4_X1 R2_SB_SB3_U445 ( .A1(R2_SB_SB3_n561), .A2(R2_SB_SB3_n560), .A3(
        R2_SB_SB3_n559), .A4(R2_SB_SB3_n558), .ZN(R2_SB_n299) );
  NAND3_X1 R2_SB_SB3_U444 ( .A1(R2_SB_SB3_n830), .A2(R2_SB_SB3_n872), .A3(
        R2_SB_SB3_n709), .ZN(R2_SB_SB3_n566) );
  NAND4_X1 R2_SB_SB3_U443 ( .A1(R2_SB_SB3_n566), .A2(R2_SB_SB3_n894), .A3(
        R2_SB_SB3_n800), .A4(R2_SB_SB3_n648), .ZN(R2_SB_SB3_n569) );
  NAND3_X1 R2_SB_SB3_U442 ( .A1(R2_SB_n305), .A2(R2_SB_n308), .A3(
        R2_SB_SB3_n744), .ZN(R2_SB_SB3_n659) );
  NAND3_X1 R2_SB_SB3_U441 ( .A1(R2_SB_SB3_n758), .A2(R2_SB_SB3_n854), .A3(
        R2_SB_SB3_n709), .ZN(R2_SB_SB3_n587) );
  NAND3_X1 R2_SB_SB3_U440 ( .A1(R2_SB_SB3_n743), .A2(R2_SB_n305), .A3(
        R2_SB_SB3_n882), .ZN(R2_SB_SB3_n592) );
  NAND4_X1 R2_SB_SB3_U439 ( .A1(R2_SB_SB3_n601), .A2(R2_SB_SB3_n600), .A3(
        R2_SB_SB3_n599), .A4(R2_SB_SB3_n598), .ZN(R2_SB_n300) );
  NAND4_X1 R2_SB_SB3_U438 ( .A1(R2_SB_SB3_n645), .A2(R2_SB_SB3_n644), .A3(
        R2_SB_SB3_n643), .A4(R2_SB_SB3_n642), .ZN(R2_SB_n301) );
  NAND3_X1 R2_SB_SB3_U437 ( .A1(R2_SB_SB3_n684), .A2(R2_SB_SB3_n843), .A3(
        R2_SB_SB3_n744), .ZN(R2_SB_SB3_n660) );
  NAND3_X1 R2_SB_SB3_U436 ( .A1(R2_SB_n305), .A2(R2_SB_SB3_n854), .A3(
        R2_SB_SB3_n792), .ZN(R2_SB_SB3_n658) );
  NAND4_X1 R2_SB_SB3_U435 ( .A1(R2_SB_SB3_n660), .A2(R2_SB_SB3_n659), .A3(
        R2_SB_SB3_n658), .A4(R2_SB_SB3_n657), .ZN(R2_SB_SB3_n668) );
  OAI33_X1 R2_SB_SB3_U434 ( .A1(R2_SB_SB3_n862), .A2(R2_SB_n312), .A3(
        R2_SB_SB3_n847), .B1(R2_SB_SB3_n903), .B2(R2_SB_SB3_n858), .B3(
        R2_SB_SB3_n830), .ZN(R2_SB_SB3_n661) );
  NAND3_X1 R2_SB_SB3_U433 ( .A1(R2_SB_SB3_n670), .A2(R2_SB_SB3_n669), .A3(
        R2_SB_SB3_n766), .ZN(R2_SB_SB3_n717) );
  NAND4_X1 R2_SB_SB3_U432 ( .A1(R2_SB_SB3_n717), .A2(R2_SB_SB3_n716), .A3(
        R2_SB_SB3_n677), .A4(R2_SB_SB3_n676), .ZN(R2_SB_SB3_n689) );
  OAI33_X1 R2_SB_SB3_U431 ( .A1(R2_SB_SB3_n839), .A2(R2_SB_SB3_n870), .A3(
        R2_SB_SB3_n883), .B1(R2_SB_SB3_n827), .B2(R2_SB_SB3_n685), .B3(
        R2_SB_SB3_n903), .ZN(R2_SB_SB3_n686) );
  NAND4_X1 R2_SB_SB3_U430 ( .A1(R2_SB_SB3_n693), .A2(R2_SB_SB3_n692), .A3(
        R2_SB_SB3_n691), .A4(R2_SB_SB3_n690), .ZN(R2_SB_n302) );
  NAND3_X1 R2_SB_SB3_U429 ( .A1(R2_SB_SB3_n845), .A2(R2_SB_SB3_n838), .A3(
        R2_SB_SB3_n829), .ZN(R2_SB_SB3_n703) );
  OAI33_X1 R2_SB_SB3_U428 ( .A1(R2_SB_SB3_n876), .A2(R2_SB_n305), .A3(
        R2_SB_SB3_n830), .B1(R2_SB_SB3_n705), .B2(R2_SB_SB3_n835), .B3(
        R2_SB_SB3_n901), .ZN(R2_SB_SB3_n706) );
  NAND3_X1 R2_SB_SB3_U427 ( .A1(R2_SB_n309), .A2(R2_SB_SB3_n714), .A3(
        R2_SB_n312), .ZN(R2_SB_SB3_n715) );
  NAND3_X1 R2_SB_SB3_U426 ( .A1(R2_SB_SB3_n717), .A2(R2_SB_SB3_n716), .A3(
        R2_SB_SB3_n715), .ZN(R2_SB_SB3_n737) );
  NAND4_X1 R2_SB_SB3_U425 ( .A1(R2_SB_SB3_n741), .A2(R2_SB_SB3_n740), .A3(
        R2_SB_SB3_n739), .A4(R2_SB_SB3_n738), .ZN(R2_SB_n303) );
  NAND3_X1 R2_SB_SB3_U424 ( .A1(R2_SB_n312), .A2(R2_SB_SB3_n854), .A3(
        R2_SB_SB3_n795), .ZN(R2_SB_SB3_n762) );
  NAND3_X1 R2_SB_SB3_U423 ( .A1(R2_SB_SB3_n763), .A2(R2_SB_SB3_n762), .A3(
        R2_SB_SB3_n761), .ZN(R2_SB_SB3_n764) );
  NAND3_X1 R2_SB_SB3_U422 ( .A1(R2_SB_n311), .A2(R2_SB_SB3_n854), .A3(
        R2_SB_SB3_n771), .ZN(R2_SB_SB3_n777) );
  NAND3_X1 R2_SB_SB3_U421 ( .A1(R2_SB_SB3_n817), .A2(R2_SB_SB3_n816), .A3(
        R2_SB_SB3_n815), .ZN(R2_SB_SB3_n820) );
  NAND4_X1 R2_SB_SB3_U420 ( .A1(R2_SB_SB3_n825), .A2(R2_SB_SB3_n824), .A3(
        R2_SB_SB3_n823), .A4(R2_SB_SB3_n822), .ZN(R2_SB_n304) );
  NOR2_X2 R2_SB_SB3_U264 ( .A1(R2_SB_SB3_n830), .A2(R2_SB_SB3_n843), .ZN(
        R2_SB_SB3_n758) );
  INV_X1 R2_SB_SB4_U466 ( .A(R2_SB_SB4_n453), .ZN(R2_SB_SB4_n452) );
  INV_X1 R2_SB_SB4_U465 ( .A(R2_SB_n290), .ZN(R2_SB_SB4_n89) );
  INV_X1 R2_SB_SB4_U419 ( .A(R2_SB_n289), .ZN(R2_SB_SB4_n453) );
  NAND2_X1 R2_SB_SB4_U418 ( .A1(R2_SB_n290), .A2(R2_SB_n295), .ZN(
        R2_SB_SB4_n705) );
  AOI22_X1 R2_SB_SB4_U417 ( .A1(R2_SB_SB4_n779), .A2(R2_SB_SB4_n760), .B1(
        R2_SB_SB4_n877), .B2(R2_SB_SB4_n792), .ZN(R2_SB_SB4_n761) );
  OAI21_X1 R2_SB_SB4_U416 ( .B1(R2_SB_SB4_n759), .B2(R2_SB_SB4_n900), .A(
        R2_SB_SB4_n758), .ZN(R2_SB_SB4_n763) );
  AOI222_X1 R2_SB_SB4_U415 ( .A1(R2_SB_SB4_n742), .A2(R2_SB_n294), .B1(
        R2_SB_SB4_n778), .B2(R2_SB_SB4_n748), .C1(R2_SB_SB4_n747), .C2(
        R2_SB_SB4_n656), .ZN(R2_SB_SB4_n657) );
  NAND2_X1 R2_SB_SB4_U414 ( .A1(R2_SB_SB4_n743), .A2(R2_SB_n296), .ZN(
        R2_SB_SB4_n472) );
  AOI21_X1 R2_SB_SB4_U413 ( .B1(R2_SB_SB4_n835), .B2(R2_SB_SB4_n837), .A(
        R2_SB_SB4_n859), .ZN(R2_SB_SB4_n474) );
  OAI21_X1 R2_SB_SB4_U412 ( .B1(R2_SB_SB4_n474), .B2(R2_SB_SB4_n473), .A(
        R2_SB_SB4_n813), .ZN(R2_SB_SB4_n475) );
  OAI22_X1 R2_SB_SB4_U411 ( .A1(R2_SB_SB4_n829), .A2(R2_SB_SB4_n847), .B1(
        R2_SB_SB4_n845), .B2(R2_SB_SB4_n826), .ZN(R2_SB_SB4_n714) );
  NOR2_X1 R2_SB_SB4_U410 ( .A1(R2_SB_n296), .A2(R2_SB_SB4_n863), .ZN(
        R2_SB_SB4_n535) );
  OAI21_X1 R2_SB_SB4_U409 ( .B1(R2_SB_SB4_n855), .B2(R2_SB_SB4_n829), .A(
        R2_SB_SB4_n745), .ZN(R2_SB_SB4_n746) );
  AOI221_X1 R2_SB_SB4_U408 ( .B1(R2_SB_SB4_n805), .B2(R2_SB_SB4_n748), .C1(
        R2_SB_SB4_n747), .C2(R2_SB_SB4_n780), .A(R2_SB_SB4_n746), .ZN(
        R2_SB_SB4_n749) );
  AOI22_X1 R2_SB_SB4_U407 ( .A1(R2_SB_SB4_n742), .A2(R2_SB_n294), .B1(
        R2_SB_SB4_n778), .B2(R2_SB_SB4_n771), .ZN(R2_SB_SB4_n750) );
  OAI211_X1 R2_SB_SB4_U406 ( .C1(R2_SB_SB4_n828), .C2(R2_SB_SB4_n847), .A(
        R2_SB_SB4_n750), .B(R2_SB_SB4_n749), .ZN(R2_SB_SB4_n751) );
  NOR2_X1 R2_SB_SB4_U405 ( .A1(R2_SB_n294), .A2(R2_SB_SB4_n830), .ZN(
        R2_SB_SB4_n724) );
  NOR2_X1 R2_SB_SB4_U404 ( .A1(R2_SB_SB4_n826), .A2(R2_SB_n292), .ZN(
        R2_SB_SB4_n463) );
  OAI22_X1 R2_SB_SB4_U403 ( .A1(R2_SB_n296), .A2(R2_SB_SB4_n876), .B1(
        R2_SB_SB4_n858), .B2(R2_SB_SB4_n901), .ZN(R2_SB_SB4_n760) );
  NOR3_X1 R2_SB_SB4_U402 ( .A1(R2_SB_SB4_n890), .A2(R2_SB_n294), .A3(
        R2_SB_n290), .ZN(R2_SB_SB4_n613) );
  OAI22_X1 R2_SB_SB4_U401 ( .A1(R2_SB_SB4_n89), .A2(R2_SB_SB4_n898), .B1(
        R2_SB_SB4_n628), .B2(R2_SB_SB4_n907), .ZN(R2_SB_SB4_n614) );
  NOR3_X1 R2_SB_SB4_U400 ( .A1(R2_SB_SB4_n614), .A2(R2_SB_SB4_n722), .A3(
        R2_SB_SB4_n613), .ZN(R2_SB_SB4_n623) );
  NOR3_X1 R2_SB_SB4_U399 ( .A1(R2_SB_SB4_n863), .A2(R2_SB_n296), .A3(
        R2_SB_SB4_n814), .ZN(R2_SB_SB4_n797) );
  AOI22_X1 R2_SB_SB4_U398 ( .A1(R2_SB_SB4_n628), .A2(R2_SB_SB4_n627), .B1(
        R2_SB_n291), .B2(R2_SB_SB4_n730), .ZN(R2_SB_SB4_n630) );
  OAI222_X1 R2_SB_SB4_U397 ( .A1(R2_SB_SB4_n837), .A2(R2_SB_SB4_n573), .B1(
        R2_SB_n289), .B2(R2_SB_SB4_n468), .C1(R2_SB_n290), .C2(R2_SB_SB4_n677), 
        .ZN(R2_SB_SB4_n483) );
  OAI221_X1 R2_SB_SB4_U396 ( .B1(R2_SB_n292), .B2(R2_SB_SB4_n581), .C1(
        R2_SB_SB4_n476), .C2(R2_SB_SB4_n878), .A(R2_SB_SB4_n475), .ZN(
        R2_SB_SB4_n482) );
  OAI22_X1 R2_SB_SB4_U395 ( .A1(R2_SB_SB4_n840), .A2(R2_SB_SB4_n800), .B1(
        R2_SB_SB4_n480), .B2(R2_SB_SB4_n453), .ZN(R2_SB_SB4_n481) );
  NOR4_X1 R2_SB_SB4_U394 ( .A1(R2_SB_SB4_n484), .A2(R2_SB_SB4_n483), .A3(
        R2_SB_SB4_n482), .A4(R2_SB_SB4_n481), .ZN(R2_SB_SB4_n485) );
  NOR2_X1 R2_SB_SB4_U393 ( .A1(R2_SB_SB4_n868), .A2(R2_SB_n296), .ZN(
        R2_SB_SB4_n680) );
  NOR2_X1 R2_SB_SB4_U392 ( .A1(R2_SB_n291), .A2(R2_SB_n293), .ZN(
        R2_SB_SB4_n646) );
  NAND2_X1 R2_SB_SB4_U391 ( .A1(R2_SB_n294), .A2(R2_SB_SB4_n872), .ZN(
        R2_SB_SB4_n770) );
  NOR2_X1 R2_SB_SB4_U390 ( .A1(R2_SB_SB4_n895), .A2(R2_SB_n292), .ZN(
        R2_SB_SB4_n783) );
  NOR2_X1 R2_SB_SB4_U389 ( .A1(R2_SB_n293), .A2(R2_SB_n294), .ZN(
        R2_SB_SB4_n617) );
  NOR2_X1 R2_SB_SB4_U388 ( .A1(R2_SB_SB4_n854), .A2(R2_SB_n291), .ZN(
        R2_SB_SB4_n811) );
  INV_X1 R2_SB_SB4_U387 ( .A(R2_SB_n296), .ZN(R2_SB_SB4_n881) );
  AOI22_X1 R2_SB_SB4_U386 ( .A1(R2_SB_n291), .A2(R2_SB_SB4_n638), .B1(
        R2_SB_SB4_n795), .B2(R2_SB_SB4_n713), .ZN(R2_SB_SB4_n711) );
  NOR2_X1 R2_SB_SB4_U385 ( .A1(R2_SB_SB4_n854), .A2(R2_SB_n294), .ZN(
        R2_SB_SB4_n694) );
  NAND2_X1 R2_SB_SB4_U384 ( .A1(R2_SB_n291), .A2(R2_SB_n294), .ZN(
        R2_SB_SB4_n608) );
  OAI221_X1 R2_SB_SB4_U383 ( .B1(R2_SB_n291), .B2(R2_SB_SB4_n551), .C1(
        R2_SB_SB4_n550), .C2(R2_SB_SB4_n910), .A(R2_SB_SB4_n902), .ZN(
        R2_SB_SB4_n552) );
  OAI221_X1 R2_SB_SB4_U382 ( .B1(R2_SB_SB4_n864), .B2(R2_SB_SB4_n838), .C1(
        R2_SB_SB4_n827), .C2(R2_SB_SB4_n849), .A(R2_SB_SB4_n615), .ZN(
        R2_SB_SB4_n553) );
  OAI221_X1 R2_SB_SB4_U381 ( .B1(R2_SB_SB4_n864), .B2(R2_SB_SB4_n835), .C1(
        R2_SB_SB4_n832), .C2(R2_SB_SB4_n853), .A(R2_SB_SB4_n546), .ZN(
        R2_SB_SB4_n554) );
  AOI221_X1 R2_SB_SB4_U380 ( .B1(R2_SB_SB4_n752), .B2(R2_SB_SB4_n554), .C1(
        R2_SB_SB4_n702), .C2(R2_SB_SB4_n553), .A(R2_SB_SB4_n552), .ZN(
        R2_SB_SB4_n559) );
  OAI22_X1 R2_SB_SB4_U379 ( .A1(R2_SB_SB4_n583), .A2(R2_SB_SB4_n826), .B1(
        R2_SB_SB4_n838), .B2(R2_SB_SB4_n891), .ZN(R2_SB_SB4_n584) );
  OAI211_X1 R2_SB_SB4_U378 ( .C1(R2_SB_SB4_n453), .C2(R2_SB_SB4_n844), .A(
        R2_SB_SB4_n835), .B(R2_SB_SB4_n847), .ZN(R2_SB_SB4_n585) );
  OAI211_X1 R2_SB_SB4_U377 ( .C1(R2_SB_n289), .C2(R2_SB_SB4_n898), .A(
        R2_SB_SB4_n582), .B(R2_SB_SB4_n581), .ZN(R2_SB_SB4_n586) );
  AOI221_X1 R2_SB_SB4_U376 ( .B1(R2_SB_n291), .B2(R2_SB_SB4_n586), .C1(
        R2_SB_SB4_n755), .C2(R2_SB_SB4_n585), .A(R2_SB_SB4_n584), .ZN(
        R2_SB_SB4_n599) );
  OAI221_X1 R2_SB_SB4_U375 ( .B1(R2_SB_SB4_n840), .B2(R2_SB_SB4_n859), .C1(
        R2_SB_SB4_n863), .C2(R2_SB_SB4_n834), .A(R2_SB_SB4_n574), .ZN(
        R2_SB_SB4_n580) );
  OAI22_X1 R2_SB_SB4_U374 ( .A1(R2_SB_n292), .A2(R2_SB_SB4_n578), .B1(
        R2_SB_SB4_n577), .B2(R2_SB_SB4_n831), .ZN(R2_SB_SB4_n579) );
  INV_X1 R2_SB_SB4_U373 ( .A(R2_SB_SB4_n573), .ZN(R2_SB_SB4_n889) );
  AOI221_X1 R2_SB_SB4_U372 ( .B1(R2_SB_SB4_n889), .B2(R2_SB_SB4_n696), .C1(
        R2_SB_SB4_n752), .C2(R2_SB_SB4_n580), .A(R2_SB_SB4_n579), .ZN(
        R2_SB_SB4_n600) );
  NOR2_X1 R2_SB_SB4_U371 ( .A1(R2_SB_n292), .A2(R2_SB_n293), .ZN(
        R2_SB_SB4_n656) );
  INV_X1 R2_SB_SB4_U370 ( .A(R2_SB_n295), .ZN(R2_SB_SB4_n872) );
  NOR3_X1 R2_SB_SB4_U369 ( .A1(R2_SB_SB4_n850), .A2(R2_SB_n293), .A3(
        R2_SB_SB4_n881), .ZN(R2_SB_SB4_n556) );
  NOR2_X1 R2_SB_SB4_U368 ( .A1(R2_SB_SB4_n830), .A2(R2_SB_n293), .ZN(
        R2_SB_SB4_n678) );
  AOI221_X1 R2_SB_SB4_U367 ( .B1(R2_SB_SB4_n806), .B2(R2_SB_SB4_n89), .C1(
        R2_SB_SB4_n805), .C2(R2_SB_SB4_n804), .A(R2_SB_SB4_n803), .ZN(
        R2_SB_SB4_n807) );
  AOI211_X1 R2_SB_SB4_U366 ( .C1(R2_SB_SB4_n799), .C2(R2_SB_SB4_n798), .A(
        R2_SB_SB4_n797), .B(R2_SB_SB4_n796), .ZN(R2_SB_SB4_n808) );
  AOI22_X1 R2_SB_SB4_U365 ( .A1(R2_SB_SB4_n793), .A2(R2_SB_SB4_n792), .B1(
        R2_SB_SB4_n791), .B2(R2_SB_SB4_n790), .ZN(R2_SB_SB4_n809) );
  OAI221_X1 R2_SB_SB4_U364 ( .B1(R2_SB_n295), .B2(R2_SB_SB4_n809), .C1(
        R2_SB_SB4_n808), .C2(R2_SB_SB4_n859), .A(R2_SB_SB4_n807), .ZN(
        R2_SB_SB4_n821) );
  NOR2_X1 R2_SB_SB4_U363 ( .A1(R2_SB_n296), .A2(R2_SB_n293), .ZN(
        R2_SB_SB4_n489) );
  OAI21_X1 R2_SB_SB4_U362 ( .B1(R2_SB_SB4_n864), .B2(R2_SB_SB4_n878), .A(
        R2_SB_SB4_n894), .ZN(R2_SB_SB4_n490) );
  AOI221_X1 R2_SB_SB4_U361 ( .B1(R2_SB_SB4_n779), .B2(R2_SB_SB4_n490), .C1(
        R2_SB_SB4_n489), .C2(R2_SB_SB4_n782), .A(R2_SB_SB4_n756), .ZN(
        R2_SB_SB4_n491) );
  AOI222_X1 R2_SB_SB4_U360 ( .A1(R2_SB_SB4_n789), .A2(R2_SB_SB4_n772), .B1(
        R2_SB_SB4_n646), .B2(R2_SB_SB4_n813), .C1(R2_SB_SB4_n709), .C2(
        R2_SB_SB4_n811), .ZN(R2_SB_SB4_n647) );
  OAI221_X1 R2_SB_SB4_U359 ( .B1(R2_SB_n290), .B2(R2_SB_SB4_n884), .C1(
        R2_SB_SB4_n453), .C2(R2_SB_SB4_n880), .A(R2_SB_SB4_n649), .ZN(
        R2_SB_SB4_n650) );
  OAI221_X1 R2_SB_SB4_U358 ( .B1(R2_SB_n292), .B2(R2_SB_SB4_n648), .C1(
        R2_SB_SB4_n845), .C2(R2_SB_SB4_n868), .A(R2_SB_SB4_n647), .ZN(
        R2_SB_SB4_n652) );
  AOI222_X1 R2_SB_SB4_U357 ( .A1(R2_SB_SB4_n781), .A2(R2_SB_SB4_n652), .B1(
        R2_SB_SB4_n651), .B2(R2_SB_SB4_n730), .C1(R2_SB_SB4_n782), .C2(
        R2_SB_SB4_n650), .ZN(R2_SB_SB4_n693) );
  NOR2_X1 R2_SB_SB4_U356 ( .A1(R2_SB_SB4_n863), .A2(R2_SB_n292), .ZN(
        R2_SB_SB4_n618) );
  NOR3_X1 R2_SB_SB4_U355 ( .A1(R2_SB_SB4_n840), .A2(R2_SB_n295), .A3(
        R2_SB_SB4_n869), .ZN(R2_SB_SB4_n575) );
  AOI221_X1 R2_SB_SB4_U354 ( .B1(R2_SB_SB4_n591), .B2(R2_SB_SB4_n453), .C1(
        R2_SB_SB4_n576), .C2(R2_SB_SB4_n684), .A(R2_SB_SB4_n575), .ZN(
        R2_SB_SB4_n578) );
  OAI211_X1 R2_SB_SB4_U353 ( .C1(R2_SB_n294), .C2(R2_SB_SB4_n848), .A(
        R2_SB_SB4_n860), .B(R2_SB_SB4_n853), .ZN(R2_SB_SB4_n662) );
  OAI21_X1 R2_SB_SB4_U352 ( .B1(R2_SB_SB4_n876), .B2(R2_SB_SB4_n853), .A(
        R2_SB_SB4_n908), .ZN(R2_SB_SB4_n663) );
  AOI221_X1 R2_SB_SB4_U351 ( .B1(R2_SB_SB4_n779), .B2(R2_SB_SB4_n663), .C1(
        R2_SB_SB4_n702), .C2(R2_SB_SB4_n662), .A(R2_SB_SB4_n661), .ZN(
        R2_SB_SB4_n664) );
  OAI222_X1 R2_SB_SB4_U350 ( .A1(R2_SB_SB4_n718), .A2(R2_SB_SB4_n907), .B1(
        R2_SB_SB4_n452), .B2(R2_SB_SB4_n664), .C1(R2_SB_SB4_n832), .C2(
        R2_SB_SB4_n802), .ZN(R2_SB_SB4_n667) );
  NOR3_X1 R2_SB_SB4_U349 ( .A1(R2_SB_SB4_n849), .A2(R2_SB_n296), .A3(
        R2_SB_SB4_n854), .ZN(R2_SB_SB4_n605) );
  OAI22_X1 R2_SB_SB4_U348 ( .A1(R2_SB_n295), .A2(R2_SB_n293), .B1(R2_SB_n294), 
        .B2(R2_SB_SB4_n883), .ZN(R2_SB_SB4_n606) );
  AOI221_X1 R2_SB_SB4_U347 ( .B1(R2_SB_SB4_n755), .B2(R2_SB_SB4_n791), .C1(
        R2_SB_SB4_n758), .C2(R2_SB_SB4_n606), .A(R2_SB_SB4_n605), .ZN(
        R2_SB_SB4_n607) );
  NOR2_X1 R2_SB_SB4_U346 ( .A1(R2_SB_SB4_n452), .A2(R2_SB_n291), .ZN(
        R2_SB_SB4_n794) );
  NOR2_X1 R2_SB_SB4_U345 ( .A1(R2_SB_n294), .A2(R2_SB_n296), .ZN(
        R2_SB_SB4_n709) );
  NOR2_X1 R2_SB_SB4_U344 ( .A1(R2_SB_SB4_n830), .A2(R2_SB_n292), .ZN(
        R2_SB_SB4_n782) );
  NOR3_X1 R2_SB_SB4_U343 ( .A1(R2_SB_SB4_n901), .A2(R2_SB_n295), .A3(
        R2_SB_SB4_n843), .ZN(R2_SB_SB4_n729) );
  AOI221_X1 R2_SB_SB4_U342 ( .B1(R2_SB_SB4_n805), .B2(R2_SB_SB4_n813), .C1(
        R2_SB_SB4_n789), .C2(R2_SB_SB4_n728), .A(R2_SB_SB4_n727), .ZN(
        R2_SB_SB4_n732) );
  AOI211_X1 R2_SB_SB4_U341 ( .C1(R2_SB_SB4_n752), .C2(R2_SB_SB4_n730), .A(
        R2_SB_SB4_n759), .B(R2_SB_SB4_n729), .ZN(R2_SB_SB4_n731) );
  OAI222_X1 R2_SB_SB4_U340 ( .A1(R2_SB_SB4_n733), .A2(R2_SB_SB4_n839), .B1(
        R2_SB_SB4_n732), .B2(R2_SB_SB4_n837), .C1(R2_SB_SB4_n731), .C2(
        R2_SB_SB4_n835), .ZN(R2_SB_SB4_n734) );
  NOR2_X1 R2_SB_SB4_U339 ( .A1(R2_SB_SB4_n854), .A2(R2_SB_n292), .ZN(
        R2_SB_SB4_n805) );
  NOR2_X1 R2_SB_SB4_U338 ( .A1(R2_SB_SB4_n872), .A2(R2_SB_n294), .ZN(
        R2_SB_SB4_n767) );
  INV_X1 R2_SB_SB4_U337 ( .A(R2_SB_n291), .ZN(R2_SB_SB4_n830) );
  NOR2_X1 R2_SB_SB4_U336 ( .A1(R2_SB_n295), .A2(R2_SB_n296), .ZN(
        R2_SB_SB4_n702) );
  NOR2_X1 R2_SB_SB4_U335 ( .A1(R2_SB_n290), .A2(R2_SB_n291), .ZN(
        R2_SB_SB4_n795) );
  NOR2_X1 R2_SB_SB4_U334 ( .A1(R2_SB_n294), .A2(R2_SB_n295), .ZN(
        R2_SB_SB4_n813) );
  NOR3_X1 R2_SB_SB4_U333 ( .A1(R2_SB_SB4_n833), .A2(R2_SB_n292), .A3(
        R2_SB_SB4_n885), .ZN(R2_SB_SB4_n639) );
  INV_X1 R2_SB_SB4_U332 ( .A(R2_SB_n293), .ZN(R2_SB_SB4_n854) );
  NOR2_X1 R2_SB_SB4_U331 ( .A1(R2_SB_SB4_n843), .A2(R2_SB_n291), .ZN(
        R2_SB_SB4_n792) );
  INV_X1 R2_SB_SB4_U330 ( .A(R2_SB_n294), .ZN(R2_SB_SB4_n863) );
  NAND2_X1 R2_SB_SB4_U329 ( .A1(R2_SB_SB4_n791), .A2(R2_SB_SB4_n772), .ZN(
        R2_SB_SB4_n775) );
  OAI21_X1 R2_SB_SB4_U328 ( .B1(R2_SB_SB4_n775), .B2(R2_SB_SB4_n774), .A(
        R2_SB_SB4_n773), .ZN(R2_SB_SB4_n776) );
  INV_X1 R2_SB_SB4_U327 ( .A(R2_SB_SB4_n776), .ZN(R2_SB_SB4_n887) );
  INV_X1 R2_SB_SB4_U326 ( .A(R2_SB_SB4_n783), .ZN(R2_SB_SB4_n897) );
  INV_X1 R2_SB_SB4_U325 ( .A(R2_SB_SB4_n678), .ZN(R2_SB_SB4_n860) );
  INV_X1 R2_SB_SB4_U324 ( .A(R2_SB_SB4_n811), .ZN(R2_SB_SB4_n855) );
  INV_X1 R2_SB_SB4_U323 ( .A(R2_SB_SB4_n463), .ZN(R2_SB_SB4_n842) );
  INV_X1 R2_SB_SB4_U322 ( .A(R2_SB_SB4_n711), .ZN(R2_SB_SB4_n909) );
  NAND2_X1 R2_SB_SB4_U321 ( .A1(R2_SB_SB4_n678), .A2(R2_SB_SB4_n781), .ZN(
        R2_SB_SB4_n615) );
  NAND2_X1 R2_SB_SB4_U320 ( .A1(R2_SB_SB4_n680), .A2(R2_SB_SB4_n810), .ZN(
        R2_SB_SB4_n581) );
  NAND2_X1 R2_SB_SB4_U319 ( .A1(R2_SB_SB4_n772), .A2(R2_SB_SB4_n684), .ZN(
        R2_SB_SB4_n785) );
  NAND2_X1 R2_SB_SB4_U318 ( .A1(R2_SB_SB4_n670), .A2(R2_SB_SB4_n881), .ZN(
        R2_SB_SB4_n773) );
  AOI22_X1 R2_SB_SB4_U317 ( .A1(R2_SB_SB4_n753), .A2(R2_SB_SB4_n771), .B1(
        R2_SB_SB4_n752), .B2(R2_SB_SB4_n751), .ZN(R2_SB_SB4_n825) );
  AOI22_X1 R2_SB_SB4_U316 ( .A1(R2_SB_n290), .A2(R2_SB_SB4_n765), .B1(
        R2_SB_SB4_n764), .B2(R2_SB_SB4_n453), .ZN(R2_SB_SB4_n824) );
  NAND2_X1 R2_SB_SB4_U315 ( .A1(R2_SB_SB4_n670), .A2(R2_SB_SB4_n872), .ZN(
        R2_SB_SB4_n801) );
  NAND2_X1 R2_SB_SB4_U314 ( .A1(R2_SB_SB4_n452), .A2(R2_SB_SB4_n843), .ZN(
        R2_SB_SB4_n548) );
  NOR2_X1 R2_SB_SB4_U313 ( .A1(R2_SB_SB4_n854), .A2(R2_SB_SB4_n827), .ZN(
        R2_SB_SB4_n793) );
  OAI21_X1 R2_SB_SB4_U312 ( .B1(R2_SB_SB4_n718), .B2(R2_SB_SB4_n588), .A(
        R2_SB_SB4_n587), .ZN(R2_SB_SB4_n597) );
  NOR4_X1 R2_SB_SB4_U311 ( .A1(R2_SB_SB4_n464), .A2(R2_SB_SB4_n886), .A3(
        R2_SB_SB4_n555), .A4(R2_SB_SB4_n639), .ZN(R2_SB_SB4_n486) );
  AOI211_X1 R2_SB_SB4_U310 ( .C1(R2_SB_SB4_n684), .C2(R2_SB_SB4_n462), .A(
        R2_SB_SB4_n461), .B(R2_SB_SB4_n460), .ZN(R2_SB_SB4_n487) );
  AOI221_X1 R2_SB_SB4_U309 ( .B1(R2_SB_SB4_n810), .B2(R2_SB_SB4_n533), .C1(
        R2_SB_SB4_n565), .C2(R2_SB_n290), .A(R2_SB_SB4_n532), .ZN(
        R2_SB_SB4_n561) );
  NOR4_X1 R2_SB_SB4_U308 ( .A1(R2_SB_SB4_n557), .A2(R2_SB_SB4_n556), .A3(
        R2_SB_SB4_n555), .A4(R2_SB_SB4_n674), .ZN(R2_SB_SB4_n558) );
  AOI221_X1 R2_SB_SB4_U307 ( .B1(R2_SB_SB4_n772), .B2(R2_SB_SB4_n572), .C1(
        R2_SB_SB4_n753), .C2(R2_SB_SB4_n758), .A(R2_SB_SB4_n571), .ZN(
        R2_SB_SB4_n601) );
  AOI211_X1 R2_SB_SB4_U306 ( .C1(R2_SB_SB4_n597), .C2(R2_SB_SB4_n453), .A(
        R2_SB_SB4_n596), .B(R2_SB_SB4_n595), .ZN(R2_SB_SB4_n598) );
  AOI221_X1 R2_SB_SB4_U305 ( .B1(R2_SB_SB4_n604), .B2(R2_SB_SB4_n877), .C1(
        R2_SB_SB4_n603), .C2(R2_SB_SB4_n679), .A(R2_SB_SB4_n602), .ZN(
        R2_SB_SB4_n645) );
  NOR4_X1 R2_SB_SB4_U304 ( .A1(R2_SB_SB4_n641), .A2(R2_SB_SB4_n640), .A3(
        R2_SB_SB4_n639), .A4(R2_SB_SB4_n673), .ZN(R2_SB_SB4_n642) );
  OAI21_X1 R2_SB_SB4_U303 ( .B1(R2_SB_SB4_n810), .B2(R2_SB_SB4_n744), .A(
        R2_SB_SB4_n743), .ZN(R2_SB_SB4_n745) );
  NOR4_X1 R2_SB_SB4_U302 ( .A1(R2_SB_SB4_n737), .A2(R2_SB_SB4_n736), .A3(
        R2_SB_SB4_n735), .A4(R2_SB_SB4_n734), .ZN(R2_SB_SB4_n738) );
  AOI211_X1 R2_SB_SB4_U301 ( .C1(R2_SB_SB4_n713), .C2(R2_SB_SB4_n758), .A(
        R2_SB_SB4_n712), .B(R2_SB_SB4_n909), .ZN(R2_SB_SB4_n739) );
  NOR4_X1 R2_SB_SB4_U300 ( .A1(R2_SB_SB4_n689), .A2(R2_SB_SB4_n688), .A3(
        R2_SB_SB4_n687), .A4(R2_SB_SB4_n686), .ZN(R2_SB_SB4_n690) );
  AOI211_X1 R2_SB_SB4_U299 ( .C1(R2_SB_SB4_n752), .C2(R2_SB_SB4_n668), .A(
        R2_SB_SB4_n667), .B(R2_SB_SB4_n666), .ZN(R2_SB_SB4_n691) );
  AOI221_X1 R2_SB_SB4_U298 ( .B1(R2_SB_SB4_n565), .B2(R2_SB_SB4_n766), .C1(
        R2_SB_SB4_n759), .C2(R2_SB_SB4_n791), .A(R2_SB_SB4_n513), .ZN(
        R2_SB_SB4_n525) );
  NOR4_X1 R2_SB_SB4_U297 ( .A1(R2_SB_SB4_n523), .A2(R2_SB_SB4_n522), .A3(
        R2_SB_SB4_n521), .A4(R2_SB_SB4_n520), .ZN(R2_SB_SB4_n524) );
  OAI221_X1 R2_SB_SB4_U296 ( .B1(R2_SB_SB4_n849), .B2(R2_SB_SB4_n770), .C1(
        R2_SB_SB4_n883), .C2(R2_SB_SB4_n608), .A(R2_SB_SB4_n567), .ZN(
        R2_SB_SB4_n568) );
  OAI21_X1 R2_SB_SB4_U295 ( .B1(R2_SB_SB4_n569), .B2(R2_SB_SB4_n568), .A(
        R2_SB_SB4_n781), .ZN(R2_SB_SB4_n570) );
  OAI21_X1 R2_SB_SB4_U294 ( .B1(R2_SB_SB4_n839), .B2(R2_SB_SB4_n892), .A(
        R2_SB_SB4_n570), .ZN(R2_SB_SB4_n571) );
  INV_X1 R2_SB_SB4_U293 ( .A(R2_SB_SB4_n780), .ZN(R2_SB_SB4_n870) );
  OAI21_X1 R2_SB_SB4_U292 ( .B1(R2_SB_SB4_n778), .B2(R2_SB_SB4_n744), .A(
        R2_SB_SB4_n696), .ZN(R2_SB_SB4_n508) );
  OAI211_X1 R2_SB_SB4_U291 ( .C1(R2_SB_SB4_n813), .C2(R2_SB_SB4_n812), .A(
        R2_SB_SB4_n811), .B(R2_SB_SB4_n810), .ZN(R2_SB_SB4_n817) );
  INV_X1 R2_SB_SB4_U290 ( .A(R2_SB_SB4_n743), .ZN(R2_SB_SB4_n851) );
  AND3_X1 R2_SB_SB4_U289 ( .A1(R2_SB_SB4_n779), .A2(R2_SB_SB4_n812), .A3(
        R2_SB_SB4_n656), .ZN(R2_SB_SB4_n87) );
  NOR3_X1 R2_SB_SB4_U288 ( .A1(R2_SB_SB4_n858), .A2(R2_SB_SB4_n665), .A3(
        R2_SB_SB4_n890), .ZN(R2_SB_SB4_n13) );
  OR3_X1 R2_SB_SB4_U287 ( .A1(R2_SB_SB4_n13), .A2(R2_SB_SB4_n675), .A3(
        R2_SB_SB4_n87), .ZN(R2_SB_SB4_n464) );
  OAI22_X1 R2_SB_SB4_U286 ( .A1(R2_SB_SB4_n872), .A2(R2_SB_SB4_n857), .B1(
        R2_SB_SB4_n854), .B2(R2_SB_SB4_n876), .ZN(R2_SB_SB4_n547) );
  INV_X1 R2_SB_SB4_U285 ( .A(R2_SB_SB4_n582), .ZN(R2_SB_SB4_n911) );
  AOI21_X1 R2_SB_SB4_U284 ( .B1(R2_SB_SB4_n781), .B2(R2_SB_SB4_n547), .A(
        R2_SB_SB4_n911), .ZN(R2_SB_SB4_n551) );
  AOI21_X1 R2_SB_SB4_U283 ( .B1(R2_SB_SB4_n754), .B2(R2_SB_SB4_n758), .A(
        R2_SB_SB4_n467), .ZN(R2_SB_SB4_n468) );
  AOI21_X1 R2_SB_SB4_U282 ( .B1(R2_SB_SB4_n778), .B2(R2_SB_SB4_n453), .A(
        R2_SB_SB4_n789), .ZN(R2_SB_SB4_n700) );
  AOI22_X1 R2_SB_SB4_U281 ( .A1(R2_SB_SB4_n725), .A2(R2_SB_SB4_n617), .B1(
        R2_SB_SB4_n766), .B2(R2_SB_SB4_n730), .ZN(R2_SB_SB4_n562) );
  AOI21_X1 R2_SB_SB4_U280 ( .B1(R2_SB_SB4_n743), .B2(R2_SB_n290), .A(
        R2_SB_SB4_n747), .ZN(R2_SB_SB4_n564) );
  OAI21_X1 R2_SB_SB4_U279 ( .B1(R2_SB_SB4_n684), .B2(R2_SB_SB4_n799), .A(
        R2_SB_SB4_n780), .ZN(R2_SB_SB4_n563) );
  OAI211_X1 R2_SB_SB4_U278 ( .C1(R2_SB_SB4_n564), .C2(R2_SB_SB4_n868), .A(
        R2_SB_SB4_n563), .B(R2_SB_SB4_n562), .ZN(R2_SB_SB4_n572) );
  OAI21_X1 R2_SB_SB4_U277 ( .B1(R2_SB_SB4_n905), .B2(R2_SB_SB4_n859), .A(
        R2_SB_SB4_n895), .ZN(R2_SB_SB4_n529) );
  AOI211_X1 R2_SB_SB4_U276 ( .C1(R2_SB_SB4_n529), .C2(R2_SB_SB4_n830), .A(
        R2_SB_SB4_n633), .B(R2_SB_SB4_n528), .ZN(R2_SB_SB4_n530) );
  AOI22_X1 R2_SB_SB4_U275 ( .A1(R2_SB_SB4_n680), .A2(R2_SB_SB4_n843), .B1(
        R2_SB_SB4_n678), .B2(R2_SB_SB4_n772), .ZN(R2_SB_SB4_n531) );
  OAI211_X1 R2_SB_SB4_U274 ( .C1(R2_SB_SB4_n905), .C2(R2_SB_SB4_n864), .A(
        R2_SB_SB4_n531), .B(R2_SB_SB4_n530), .ZN(R2_SB_SB4_n533) );
  OAI21_X1 R2_SB_SB4_U273 ( .B1(R2_SB_SB4_n755), .B2(R2_SB_SB4_n754), .A(
        R2_SB_SB4_n782), .ZN(R2_SB_SB4_n757) );
  INV_X1 R2_SB_SB4_U272 ( .A(R2_SB_SB4_n756), .ZN(R2_SB_SB4_n899) );
  OAI211_X1 R2_SB_SB4_U271 ( .C1(R2_SB_SB4_n845), .C2(R2_SB_SB4_n880), .A(
        R2_SB_SB4_n757), .B(R2_SB_SB4_n899), .ZN(R2_SB_SB4_n765) );
  INV_X1 R2_SB_SB4_U270 ( .A(R2_SB_SB4_n696), .ZN(R2_SB_SB4_n836) );
  AOI21_X1 R2_SB_SB4_U269 ( .B1(R2_SB_SB4_n843), .B2(R2_SB_SB4_n835), .A(
        R2_SB_SB4_n879), .ZN(R2_SB_SB4_n595) );
  NAND2_X1 R2_SB_SB4_U268 ( .A1(R2_SB_SB4_n634), .A2(R2_SB_SB4_n805), .ZN(
        R2_SB_SB4_n800) );
  NAND2_X1 R2_SB_SB4_U267 ( .A1(R2_SB_SB4_n772), .A2(R2_SB_SB4_n507), .ZN(
        R2_SB_SB4_n648) );
  AOI21_X1 R2_SB_SB4_U266 ( .B1(R2_SB_SB4_n849), .B2(R2_SB_SB4_n608), .A(
        R2_SB_SB4_n878), .ZN(R2_SB_SB4_n528) );
  INV_X1 R2_SB_SB4_U265 ( .A(R2_SB_SB4_n794), .ZN(R2_SB_SB4_n837) );
  NOR2_X1 R2_SB_SB4_U263 ( .A1(R2_SB_SB4_n770), .A2(R2_SB_SB4_n833), .ZN(
        R2_SB_SB4_n651) );
  INV_X1 R2_SB_SB4_U262 ( .A(R2_SB_SB4_n798), .ZN(R2_SB_SB4_n901) );
  INV_X1 R2_SB_SB4_U261 ( .A(R2_SB_SB4_n813), .ZN(R2_SB_SB4_n876) );
  AOI22_X1 R2_SB_SB4_U260 ( .A1(R2_SB_SB4_n696), .A2(R2_SB_SB4_n789), .B1(
        R2_SB_SB4_n778), .B2(R2_SB_SB4_n779), .ZN(R2_SB_SB4_n612) );
  AOI22_X1 R2_SB_SB4_U259 ( .A1(R2_SB_SB4_n795), .A2(R2_SB_SB4_n798), .B1(
        R2_SB_SB4_n767), .B2(R2_SB_SB4_n766), .ZN(R2_SB_SB4_n768) );
  NAND2_X1 R2_SB_SB4_U258 ( .A1(R2_SB_SB4_n865), .A2(R2_SB_SB4_n853), .ZN(
        R2_SB_SB4_n495) );
  AOI22_X1 R2_SB_SB4_U257 ( .A1(R2_SB_SB4_n684), .A2(R2_SB_SB4_n495), .B1(
        R2_SB_SB4_n696), .B2(R2_SB_SB4_n618), .ZN(R2_SB_SB4_n496) );
  INV_X1 R2_SB_SB4_U256 ( .A(R2_SB_SB4_n805), .ZN(R2_SB_SB4_n857) );
  NAND2_X1 R2_SB_SB4_U255 ( .A1(R2_SB_SB4_n843), .A2(R2_SB_SB4_n863), .ZN(
        R2_SB_SB4_n774) );
  AOI22_X1 R2_SB_SB4_U254 ( .A1(R2_SB_SB4_n798), .A2(R2_SB_SB4_n627), .B1(
        R2_SB_SB4_n743), .B2(R2_SB_SB4_n752), .ZN(R2_SB_SB4_n567) );
  INV_X1 R2_SB_SB4_U253 ( .A(R2_SB_SB4_n767), .ZN(R2_SB_SB4_n874) );
  NOR2_X1 R2_SB_SB4_U252 ( .A1(R2_SB_SB4_n795), .A2(R2_SB_SB4_n794), .ZN(
        R2_SB_SB4_n814) );
  INV_X1 R2_SB_SB4_U251 ( .A(R2_SB_SB4_n694), .ZN(R2_SB_SB4_n869) );
  NOR2_X1 R2_SB_SB4_U250 ( .A1(R2_SB_SB4_n830), .A2(R2_SB_SB4_n684), .ZN(
        R2_SB_SB4_n665) );
  NOR2_X1 R2_SB_SB4_U249 ( .A1(R2_SB_SB4_n843), .A2(R2_SB_n290), .ZN(
        R2_SB_SB4_n604) );
  NOR2_X1 R2_SB_SB4_U248 ( .A1(R2_SB_SB4_n863), .A2(R2_SB_SB4_n858), .ZN(
        R2_SB_SB4_n790) );
  NAND2_X1 R2_SB_SB4_U247 ( .A1(R2_SB_SB4_n752), .A2(R2_SB_SB4_n507), .ZN(
        R2_SB_SB4_n802) );
  AOI21_X1 R2_SB_SB4_U246 ( .B1(R2_SB_SB4_n789), .B2(R2_SB_SB4_n798), .A(
        R2_SB_SB4_n783), .ZN(R2_SB_SB4_n721) );
  OAI21_X1 R2_SB_SB4_U245 ( .B1(R2_SB_SB4_n747), .B2(R2_SB_SB4_n843), .A(
        R2_SB_SB4_n759), .ZN(R2_SB_SB4_n719) );
  OR3_X1 R2_SB_SB4_U244 ( .A1(R2_SB_SB4_n718), .A2(R2_SB_SB4_n452), .A3(
        R2_SB_SB4_n802), .ZN(R2_SB_SB4_n720) );
  OAI211_X1 R2_SB_SB4_U243 ( .C1(R2_SB_SB4_n721), .C2(R2_SB_SB4_n826), .A(
        R2_SB_SB4_n720), .B(R2_SB_SB4_n719), .ZN(R2_SB_SB4_n736) );
  AOI22_X1 R2_SB_SB4_U242 ( .A1(R2_SB_SB4_n678), .A2(R2_SB_SB4_n767), .B1(
        R2_SB_SB4_n900), .B2(R2_SB_SB4_n843), .ZN(R2_SB_SB4_n683) );
  OAI21_X1 R2_SB_SB4_U241 ( .B1(R2_SB_SB4_n794), .B2(R2_SB_SB4_n791), .A(
        R2_SB_SB4_n882), .ZN(R2_SB_SB4_n681) );
  OAI21_X1 R2_SB_SB4_U240 ( .B1(R2_SB_SB4_n680), .B2(R2_SB_SB4_n679), .A(
        R2_SB_SB4_n696), .ZN(R2_SB_SB4_n682) );
  OAI211_X1 R2_SB_SB4_U239 ( .C1(R2_SB_SB4_n683), .C2(R2_SB_SB4_n829), .A(
        R2_SB_SB4_n682), .B(R2_SB_SB4_n681), .ZN(R2_SB_SB4_n688) );
  NOR3_X1 R2_SB_SB4_U238 ( .A1(R2_SB_SB4_n848), .A2(R2_SB_SB4_n452), .A3(
        R2_SB_SB4_n863), .ZN(R2_SB_SB4_n540) );
  OAI22_X1 R2_SB_SB4_U237 ( .A1(R2_SB_SB4_n858), .A2(R2_SB_SB4_n838), .B1(
        R2_SB_SB4_n857), .B2(R2_SB_SB4_n840), .ZN(R2_SB_SB4_n541) );
  AOI21_X1 R2_SB_SB4_U236 ( .B1(R2_SB_n290), .B2(R2_SB_SB4_n548), .A(
        R2_SB_SB4_n862), .ZN(R2_SB_SB4_n539) );
  NOR3_X1 R2_SB_SB4_U235 ( .A1(R2_SB_SB4_n541), .A2(R2_SB_SB4_n540), .A3(
        R2_SB_SB4_n539), .ZN(R2_SB_SB4_n542) );
  AOI21_X1 R2_SB_SB4_U234 ( .B1(R2_SB_SB4_n730), .B2(R2_SB_SB4_n709), .A(
        R2_SB_SB4_n753), .ZN(R2_SB_SB4_n733) );
  INV_X1 R2_SB_SB4_U233 ( .A(R2_SB_SB4_n791), .ZN(R2_SB_SB4_n840) );
  NOR3_X1 R2_SB_SB4_U232 ( .A1(R2_SB_SB4_n828), .A2(R2_SB_SB4_n856), .A3(
        R2_SB_SB4_n876), .ZN(R2_SB_SB4_n819) );
  AOI21_X1 R2_SB_SB4_U231 ( .B1(R2_SB_SB4_n845), .B2(R2_SB_SB4_n837), .A(
        R2_SB_SB4_n906), .ZN(R2_SB_SB4_n818) );
  NOR4_X1 R2_SB_SB4_U230 ( .A1(R2_SB_SB4_n821), .A2(R2_SB_SB4_n820), .A3(
        R2_SB_SB4_n819), .A4(R2_SB_SB4_n818), .ZN(R2_SB_SB4_n822) );
  INV_X1 R2_SB_SB4_U229 ( .A(R2_SB_SB4_n789), .ZN(R2_SB_SB4_n853) );
  NOR2_X1 R2_SB_SB4_U228 ( .A1(R2_SB_SB4_n743), .A2(R2_SB_SB4_n603), .ZN(
        R2_SB_SB4_n718) );
  AOI221_X1 R2_SB_SB4_U227 ( .B1(R2_SB_SB4_n877), .B2(R2_SB_SB4_n684), .C1(
        R2_SB_SB4_n591), .C2(R2_SB_SB4_n89), .A(R2_SB_SB4_n590), .ZN(
        R2_SB_SB4_n593) );
  AOI22_X1 R2_SB_SB4_U226 ( .A1(R2_SB_SB4_n810), .A2(R2_SB_SB4_n589), .B1(
        R2_SB_SB4_n798), .B2(R2_SB_SB4_n723), .ZN(R2_SB_SB4_n594) );
  OAI221_X1 R2_SB_SB4_U225 ( .B1(R2_SB_SB4_n594), .B2(R2_SB_SB4_n859), .C1(
        R2_SB_SB4_n593), .C2(R2_SB_SB4_n849), .A(R2_SB_SB4_n592), .ZN(
        R2_SB_SB4_n596) );
  INV_X1 R2_SB_SB4_U224 ( .A(R2_SB_SB4_n744), .ZN(R2_SB_SB4_n868) );
  OAI21_X1 R2_SB_SB4_U223 ( .B1(R2_SB_SB4_n779), .B2(R2_SB_SB4_n453), .A(
        R2_SB_SB4_n656), .ZN(R2_SB_SB4_n503) );
  NOR2_X1 R2_SB_SB4_U222 ( .A1(R2_SB_SB4_n618), .A2(R2_SB_SB4_n780), .ZN(
        R2_SB_SB4_n504) );
  OAI221_X1 R2_SB_SB4_U221 ( .B1(R2_SB_SB4_n504), .B2(R2_SB_SB4_n840), .C1(
        R2_SB_SB4_n869), .C2(R2_SB_SB4_n852), .A(R2_SB_SB4_n503), .ZN(
        R2_SB_SB4_n505) );
  INV_X1 R2_SB_SB4_U220 ( .A(R2_SB_SB4_n617), .ZN(R2_SB_SB4_n862) );
  AOI21_X1 R2_SB_SB4_U219 ( .B1(R2_SB_SB4_n828), .B2(R2_SB_SB4_n850), .A(
        R2_SB_SB4_n879), .ZN(R2_SB_SB4_n459) );
  AOI221_X1 R2_SB_SB4_U218 ( .B1(R2_SB_SB4_n463), .B2(R2_SB_SB4_n591), .C1(
        R2_SB_SB4_n514), .C2(R2_SB_SB4_n766), .A(R2_SB_SB4_n459), .ZN(
        R2_SB_SB4_n488) );
  OAI222_X1 R2_SB_SB4_U217 ( .A1(R2_SB_SB4_n623), .A2(R2_SB_SB4_n851), .B1(
        R2_SB_SB4_n622), .B2(R2_SB_SB4_n883), .C1(R2_SB_SB4_n621), .C2(
        R2_SB_SB4_n905), .ZN(R2_SB_SB4_n624) );
  OAI221_X1 R2_SB_SB4_U216 ( .B1(R2_SB_SB4_n903), .B2(R2_SB_SB4_n844), .C1(
        R2_SB_SB4_n848), .C2(R2_SB_SB4_n910), .A(R2_SB_SB4_n607), .ZN(
        R2_SB_SB4_n626) );
  OAI211_X1 R2_SB_SB4_U215 ( .C1(R2_SB_SB4_n857), .C2(R2_SB_SB4_n831), .A(
        R2_SB_SB4_n612), .B(R2_SB_SB4_n611), .ZN(R2_SB_SB4_n625) );
  AOI221_X1 R2_SB_SB4_U214 ( .B1(R2_SB_SB4_n452), .B2(R2_SB_SB4_n626), .C1(
        R2_SB_SB4_n752), .C2(R2_SB_SB4_n625), .A(R2_SB_SB4_n624), .ZN(
        R2_SB_SB4_n644) );
  OAI22_X1 R2_SB_SB4_U213 ( .A1(R2_SB_SB4_n733), .A2(R2_SB_SB4_n837), .B1(
        R2_SB_SB4_n842), .B2(R2_SB_SB4_n884), .ZN(R2_SB_SB4_n653) );
  OAI22_X1 R2_SB_SB4_U212 ( .A1(R2_SB_SB4_n858), .A2(R2_SB_SB4_n834), .B1(
        R2_SB_n290), .B2(R2_SB_SB4_n859), .ZN(R2_SB_SB4_n654) );
  OAI21_X1 R2_SB_SB4_U211 ( .B1(R2_SB_SB4_n903), .B2(R2_SB_SB4_n859), .A(
        R2_SB_SB4_n895), .ZN(R2_SB_SB4_n655) );
  AOI221_X1 R2_SB_SB4_U210 ( .B1(R2_SB_SB4_n795), .B2(R2_SB_SB4_n655), .C1(
        R2_SB_SB4_n702), .C2(R2_SB_SB4_n654), .A(R2_SB_SB4_n653), .ZN(
        R2_SB_SB4_n692) );
  AOI221_X1 R2_SB_SB4_U209 ( .B1(R2_SB_SB4_n684), .B2(R2_SB_SB4_n536), .C1(
        R2_SB_SB4_n535), .C2(R2_SB_SB4_n628), .A(R2_SB_SB4_n534), .ZN(
        R2_SB_SB4_n537) );
  OAI222_X1 R2_SB_SB4_U208 ( .A1(R2_SB_SB4_n543), .A2(R2_SB_SB4_n847), .B1(
        R2_SB_SB4_n835), .B2(R2_SB_SB4_n573), .C1(R2_SB_SB4_n542), .C2(
        R2_SB_SB4_n883), .ZN(R2_SB_SB4_n544) );
  OAI221_X1 R2_SB_SB4_U207 ( .B1(R2_SB_SB4_n89), .B2(R2_SB_SB4_n588), .C1(
        R2_SB_n289), .C2(R2_SB_SB4_n910), .A(R2_SB_SB4_n537), .ZN(
        R2_SB_SB4_n545) );
  AOI221_X1 R2_SB_SB4_U206 ( .B1(R2_SB_SB4_n792), .B2(R2_SB_SB4_n545), .C1(
        R2_SB_SB4_n753), .C2(R2_SB_SB4_n791), .A(R2_SB_SB4_n544), .ZN(
        R2_SB_SB4_n560) );
  AOI22_X1 R2_SB_SB4_U205 ( .A1(R2_SB_SB4_n798), .A2(R2_SB_SB4_n708), .B1(
        R2_SB_SB4_n795), .B2(R2_SB_SB4_n767), .ZN(R2_SB_SB4_n631) );
  AOI21_X1 R2_SB_SB4_U204 ( .B1(R2_SB_SB4_n755), .B2(R2_SB_SB4_n758), .A(
        R2_SB_SB4_n756), .ZN(R2_SB_SB4_n629) );
  OAI222_X1 R2_SB_SB4_U203 ( .A1(R2_SB_SB4_n631), .A2(R2_SB_SB4_n857), .B1(
        R2_SB_SB4_n630), .B2(R2_SB_SB4_n875), .C1(R2_SB_n290), .C2(
        R2_SB_SB4_n629), .ZN(R2_SB_SB4_n632) );
  AOI221_X1 R2_SB_SB4_U202 ( .B1(R2_SB_SB4_n725), .B2(R2_SB_SB4_n728), .C1(
        R2_SB_SB4_n651), .C2(R2_SB_SB4_n789), .A(R2_SB_SB4_n632), .ZN(
        R2_SB_SB4_n643) );
  OAI222_X1 R2_SB_SB4_U201 ( .A1(R2_SB_SB4_n865), .A2(R2_SB_SB4_n785), .B1(
        R2_SB_SB4_n784), .B2(R2_SB_SB4_n905), .C1(R2_SB_SB4_n827), .C2(
        R2_SB_SB4_n897), .ZN(R2_SB_SB4_n786) );
  OAI211_X1 R2_SB_SB4_U200 ( .C1(R2_SB_SB4_n829), .C2(R2_SB_SB4_n770), .A(
        R2_SB_SB4_n769), .B(R2_SB_SB4_n768), .ZN(R2_SB_SB4_n788) );
  OAI211_X1 R2_SB_SB4_U199 ( .C1(R2_SB_SB4_n895), .C2(R2_SB_SB4_n848), .A(
        R2_SB_SB4_n777), .B(R2_SB_SB4_n887), .ZN(R2_SB_SB4_n787) );
  AOI221_X1 R2_SB_SB4_U198 ( .B1(R2_SB_SB4_n789), .B2(R2_SB_SB4_n788), .C1(
        R2_SB_n289), .C2(R2_SB_SB4_n787), .A(R2_SB_SB4_n786), .ZN(
        R2_SB_SB4_n823) );
  INV_X1 R2_SB_SB4_U197 ( .A(R2_SB_SB4_n656), .ZN(R2_SB_SB4_n859) );
  AOI211_X1 R2_SB_SB4_U196 ( .C1(R2_SB_SB4_n789), .C2(R2_SB_SB4_n812), .A(
        R2_SB_SB4_n882), .B(R2_SB_SB4_n727), .ZN(R2_SB_SB4_n577) );
  AOI211_X1 R2_SB_SB4_U195 ( .C1(R2_SB_SB4_n744), .C2(R2_SB_SB4_n843), .A(
        R2_SB_SB4_n730), .B(R2_SB_SB4_n792), .ZN(R2_SB_SB4_n509) );
  AOI21_X1 R2_SB_SB4_U194 ( .B1(R2_SB_SB4_n854), .B2(R2_SB_SB4_n881), .A(
        R2_SB_SB4_n767), .ZN(R2_SB_SB4_n477) );
  OAI222_X1 R2_SB_SB4_U193 ( .A1(R2_SB_SB4_n843), .A2(R2_SB_SB4_n885), .B1(
        R2_SB_SB4_n477), .B2(R2_SB_SB4_n845), .C1(R2_SB_SB4_n864), .C2(
        R2_SB_SB4_n878), .ZN(R2_SB_SB4_n479) );
  OAI22_X1 R2_SB_SB4_U192 ( .A1(R2_SB_SB4_n849), .A2(R2_SB_SB4_n648), .B1(
        R2_SB_SB4_n862), .B2(R2_SB_SB4_n844), .ZN(R2_SB_SB4_n478) );
  AOI211_X1 R2_SB_SB4_U191 ( .C1(R2_SB_SB4_n791), .C2(R2_SB_SB4_n812), .A(
        R2_SB_SB4_n479), .B(R2_SB_SB4_n478), .ZN(R2_SB_SB4_n480) );
  NOR3_X1 R2_SB_SB4_U190 ( .A1(R2_SB_SB4_n838), .A2(R2_SB_n289), .A3(
        R2_SB_SB4_n864), .ZN(R2_SB_SB4_n610) );
  AOI21_X1 R2_SB_SB4_U189 ( .B1(R2_SB_SB4_n858), .B2(R2_SB_SB4_n608), .A(
        R2_SB_SB4_n827), .ZN(R2_SB_SB4_n609) );
  AOI211_X1 R2_SB_SB4_U188 ( .C1(R2_SB_SB4_n646), .C2(R2_SB_SB4_n781), .A(
        R2_SB_SB4_n610), .B(R2_SB_SB4_n609), .ZN(R2_SB_SB4_n611) );
  INV_X1 R2_SB_SB4_U187 ( .A(R2_SB_SB4_n752), .ZN(R2_SB_SB4_n878) );
  NOR2_X1 R2_SB_SB4_U186 ( .A1(R2_SB_SB4_n857), .A2(R2_SB_SB4_n863), .ZN(
        R2_SB_SB4_n670) );
  INV_X1 R2_SB_SB4_U185 ( .A(R2_SB_SB4_n772), .ZN(R2_SB_SB4_n883) );
  INV_X1 R2_SB_SB4_U184 ( .A(R2_SB_SB4_n618), .ZN(R2_SB_SB4_n864) );
  OAI21_X1 R2_SB_SB4_U183 ( .B1(R2_SB_SB4_n856), .B2(R2_SB_SB4_n874), .A(
        R2_SB_SB4_n893), .ZN(R2_SB_SB4_n516) );
  AOI21_X1 R2_SB_SB4_U182 ( .B1(R2_SB_SB4_n781), .B2(R2_SB_SB4_n516), .A(
        R2_SB_SB4_n515), .ZN(R2_SB_SB4_n517) );
  AOI21_X1 R2_SB_SB4_U181 ( .B1(R2_SB_SB4_n900), .B2(R2_SB_SB4_n603), .A(
        R2_SB_SB4_n783), .ZN(R2_SB_SB4_n518) );
  OAI221_X1 R2_SB_SB4_U180 ( .B1(R2_SB_SB4_n518), .B2(R2_SB_SB4_n453), .C1(
        R2_SB_SB4_n838), .C2(R2_SB_SB4_n904), .A(R2_SB_SB4_n517), .ZN(
        R2_SB_SB4_n523) );
  AOI21_X1 R2_SB_SB4_U179 ( .B1(R2_SB_SB4_n646), .B2(R2_SB_SB4_n634), .A(
        R2_SB_SB4_n633), .ZN(R2_SB_SB4_n636) );
  OAI21_X1 R2_SB_SB4_U178 ( .B1(R2_SB_SB4_n747), .B2(R2_SB_SB4_n799), .A(
        R2_SB_SB4_n882), .ZN(R2_SB_SB4_n635) );
  NAND2_X1 R2_SB_SB4_U177 ( .A1(R2_SB_SB4_n828), .A2(R2_SB_SB4_n843), .ZN(
        R2_SB_SB4_n637) );
  OAI221_X1 R2_SB_SB4_U176 ( .B1(R2_SB_SB4_n910), .B2(R2_SB_SB4_n637), .C1(
        R2_SB_SB4_n636), .C2(R2_SB_SB4_n829), .A(R2_SB_SB4_n635), .ZN(
        R2_SB_SB4_n641) );
  OAI22_X1 R2_SB_SB4_U175 ( .A1(R2_SB_SB4_n857), .A2(R2_SB_SB4_n838), .B1(
        R2_SB_SB4_n832), .B2(R2_SB_SB4_n865), .ZN(R2_SB_SB4_n469) );
  OAI21_X1 R2_SB_SB4_U174 ( .B1(R2_SB_n290), .B2(R2_SB_SB4_n845), .A(
        R2_SB_SB4_n849), .ZN(R2_SB_SB4_n471) );
  AOI221_X1 R2_SB_SB4_U173 ( .B1(R2_SB_SB4_n744), .B2(R2_SB_SB4_n471), .C1(
        R2_SB_SB4_n470), .C2(R2_SB_SB4_n863), .A(R2_SB_SB4_n469), .ZN(
        R2_SB_SB4_n476) );
  AOI221_X1 R2_SB_SB4_U172 ( .B1(R2_SB_SB4_n882), .B2(R2_SB_SB4_n792), .C1(
        R2_SB_SB4_n627), .C2(R2_SB_SB4_n702), .A(R2_SB_SB4_n698), .ZN(
        R2_SB_SB4_n583) );
  NOR2_X1 R2_SB_SB4_U171 ( .A1(R2_SB_SB4_n813), .A2(R2_SB_SB4_n694), .ZN(
        R2_SB_SB4_n695) );
  OAI221_X1 R2_SB_SB4_U170 ( .B1(R2_SB_SB4_n695), .B2(R2_SB_SB4_n851), .C1(
        R2_SB_SB4_n856), .C2(R2_SB_SB4_n878), .A(R2_SB_SB4_n904), .ZN(
        R2_SB_SB4_n697) );
  INV_X1 R2_SB_SB4_U169 ( .A(R2_SB_SB4_n801), .ZN(R2_SB_SB4_n873) );
  AOI222_X1 R2_SB_SB4_U168 ( .A1(R2_SB_SB4_n771), .A2(R2_SB_SB4_n698), .B1(
        R2_SB_SB4_n781), .B2(R2_SB_SB4_n697), .C1(R2_SB_SB4_n696), .C2(
        R2_SB_SB4_n873), .ZN(R2_SB_SB4_n741) );
  AOI22_X1 R2_SB_SB4_U167 ( .A1(R2_SB_SB4_n758), .A2(R2_SB_SB4_n694), .B1(
        R2_SB_SB4_n779), .B2(R2_SB_SB4_n863), .ZN(R2_SB_SB4_n619) );
  OAI222_X1 R2_SB_SB4_U166 ( .A1(R2_SB_SB4_n864), .A2(R2_SB_SB4_n833), .B1(
        R2_SB_n289), .B2(R2_SB_SB4_n619), .C1(R2_SB_SB4_n858), .C2(
        R2_SB_SB4_n839), .ZN(R2_SB_SB4_n620) );
  AOI221_X1 R2_SB_SB4_U165 ( .B1(R2_SB_SB4_n789), .B2(R2_SB_SB4_n628), .C1(
        R2_SB_SB4_n778), .C2(R2_SB_SB4_n771), .A(R2_SB_SB4_n620), .ZN(
        R2_SB_SB4_n621) );
  NAND2_X1 R2_SB_SB4_U164 ( .A1(R2_SB_SB4_n848), .A2(R2_SB_SB4_n841), .ZN(
        R2_SB_SB4_n616) );
  INV_X1 R2_SB_SB4_U163 ( .A(R2_SB_SB4_n615), .ZN(R2_SB_SB4_n861) );
  AOI221_X1 R2_SB_SB4_U162 ( .B1(R2_SB_SB4_n747), .B2(R2_SB_SB4_n618), .C1(
        R2_SB_SB4_n617), .C2(R2_SB_SB4_n616), .A(R2_SB_SB4_n861), .ZN(
        R2_SB_SB4_n622) );
  OAI221_X1 R2_SB_SB4_U161 ( .B1(R2_SB_SB4_n870), .B2(R2_SB_SB4_n838), .C1(
        R2_SB_SB4_n840), .C2(R2_SB_SB4_n868), .A(R2_SB_SB4_n496), .ZN(
        R2_SB_SB4_n497) );
  OAI211_X1 R2_SB_SB4_U160 ( .C1(R2_SB_SB4_n879), .C2(R2_SB_SB4_n844), .A(
        R2_SB_SB4_n711), .B(R2_SB_SB4_n491), .ZN(R2_SB_SB4_n499) );
  AOI222_X1 R2_SB_SB4_U159 ( .A1(R2_SB_SB4_n499), .A2(R2_SB_SB4_n453), .B1(
        R2_SB_SB4_n498), .B2(R2_SB_SB4_n854), .C1(R2_SB_SB4_n752), .C2(
        R2_SB_SB4_n497), .ZN(R2_SB_SB4_n527) );
  OAI222_X1 R2_SB_SB4_U158 ( .A1(R2_SB_SB4_n865), .A2(R2_SB_SB4_n838), .B1(
        R2_SB_SB4_n699), .B2(R2_SB_SB4_n868), .C1(R2_SB_n290), .C2(
        R2_SB_SB4_n858), .ZN(R2_SB_SB4_n704) );
  OAI22_X1 R2_SB_SB4_U157 ( .A1(R2_SB_SB4_n864), .A2(R2_SB_SB4_n839), .B1(
        R2_SB_SB4_n700), .B2(R2_SB_SB4_n833), .ZN(R2_SB_SB4_n701) );
  AOI222_X1 R2_SB_SB4_U156 ( .A1(R2_SB_SB4_n772), .A2(R2_SB_SB4_n704), .B1(
        R2_SB_SB4_n882), .B2(R2_SB_SB4_n703), .C1(R2_SB_SB4_n702), .C2(
        R2_SB_SB4_n701), .ZN(R2_SB_SB4_n740) );
  NOR2_X1 R2_SB_SB4_U155 ( .A1(R2_SB_SB4_n881), .A2(R2_SB_SB4_n863), .ZN(
        R2_SB_SB4_n634) );
  OAI222_X1 R2_SB_SB4_U154 ( .A1(R2_SB_n290), .A2(R2_SB_SB4_n875), .B1(
        R2_SB_SB4_n883), .B2(R2_SB_SB4_n826), .C1(R2_SB_SB4_n905), .C2(
        R2_SB_SB4_n831), .ZN(R2_SB_SB4_n707) );
  AOI211_X1 R2_SB_SB4_U153 ( .C1(R2_SB_SB4_n709), .C2(R2_SB_SB4_n708), .A(
        R2_SB_SB4_n707), .B(R2_SB_SB4_n706), .ZN(R2_SB_SB4_n710) );
  OAI222_X1 R2_SB_SB4_U152 ( .A1(R2_SB_SB4_n833), .A2(R2_SB_SB4_n898), .B1(
        R2_SB_SB4_n710), .B2(R2_SB_SB4_n859), .C1(R2_SB_SB4_n832), .C2(
        R2_SB_SB4_n800), .ZN(R2_SB_SB4_n712) );
  INV_X1 R2_SB_SB4_U151 ( .A(R2_SB_SB4_n792), .ZN(R2_SB_SB4_n845) );
  OAI221_X1 R2_SB_SB4_U150 ( .B1(R2_SB_SB4_n833), .B2(R2_SB_SB4_n774), .C1(
        R2_SB_SB4_n509), .C2(R2_SB_SB4_n829), .A(R2_SB_SB4_n508), .ZN(
        R2_SB_SB4_n510) );
  AOI221_X1 R2_SB_SB4_U149 ( .B1(R2_SB_SB4_n507), .B2(R2_SB_SB4_n506), .C1(
        R2_SB_SB4_n780), .C2(R2_SB_SB4_n684), .A(R2_SB_SB4_n505), .ZN(
        R2_SB_SB4_n512) );
  AOI221_X1 R2_SB_SB4_U148 ( .B1(R2_SB_SB4_n743), .B2(R2_SB_SB4_n684), .C1(
        R2_SB_SB4_n780), .C2(R2_SB_SB4_n627), .A(R2_SB_SB4_n510), .ZN(
        R2_SB_SB4_n511) );
  OAI222_X1 R2_SB_SB4_U147 ( .A1(R2_SB_SB4_n512), .A2(R2_SB_SB4_n905), .B1(
        R2_SB_SB4_n511), .B2(R2_SB_SB4_n883), .C1(R2_SB_SB4_n884), .C2(
        R2_SB_SB4_n844), .ZN(R2_SB_SB4_n513) );
  INV_X1 R2_SB_SB4_U146 ( .A(R2_SB_SB4_n659), .ZN(R2_SB_SB4_n867) );
  AOI221_X1 R2_SB_SB4_U145 ( .B1(R2_SB_SB4_n794), .B2(R2_SB_SB4_n730), .C1(
        R2_SB_SB4_n742), .C2(R2_SB_SB4_n780), .A(R2_SB_SB4_n867), .ZN(
        R2_SB_SB4_n574) );
  NOR4_X1 R2_SB_SB4_U144 ( .A1(R2_SB_SB4_n452), .A2(R2_SB_SB4_n872), .A3(
        R2_SB_SB4_n849), .A4(R2_SB_SB4_n862), .ZN(R2_SB_SB4_n640) );
  NOR2_X1 R2_SB_SB4_U143 ( .A1(R2_SB_SB4_n89), .A2(R2_SB_SB4_n843), .ZN(
        R2_SB_SB4_n603) );
  NOR2_X1 R2_SB_SB4_U142 ( .A1(R2_SB_SB4_n872), .A2(R2_SB_SB4_n863), .ZN(
        R2_SB_SB4_n812) );
  NOR2_X1 R2_SB_SB4_U141 ( .A1(R2_SB_SB4_n863), .A2(R2_SB_SB4_n854), .ZN(
        R2_SB_SB4_n507) );
  AOI222_X1 R2_SB_SB4_U140 ( .A1(R2_SB_SB4_n782), .A2(R2_SB_SB4_n781), .B1(
        R2_SB_SB4_n780), .B2(R2_SB_SB4_n779), .C1(R2_SB_SB4_n778), .C2(
        R2_SB_SB4_n791), .ZN(R2_SB_SB4_n784) );
  INV_X1 R2_SB_SB4_U139 ( .A(R2_SB_SB4_n795), .ZN(R2_SB_SB4_n838) );
  AOI22_X1 R2_SB_SB4_U138 ( .A1(R2_SB_SB4_n724), .A2(R2_SB_SB4_n810), .B1(
        R2_SB_SB4_n744), .B2(R2_SB_SB4_n723), .ZN(R2_SB_SB4_n726) );
  INV_X1 R2_SB_SB4_U137 ( .A(R2_SB_SB4_n722), .ZN(R2_SB_SB4_n896) );
  INV_X1 R2_SB_SB4_U136 ( .A(R2_SB_SB4_n725), .ZN(R2_SB_SB4_n846) );
  OAI222_X1 R2_SB_SB4_U135 ( .A1(R2_SB_SB4_n849), .A2(R2_SB_SB4_n896), .B1(
        R2_SB_SB4_n726), .B2(R2_SB_SB4_n878), .C1(R2_SB_SB4_n846), .C2(
        R2_SB_SB4_n910), .ZN(R2_SB_SB4_n735) );
  OAI222_X1 R2_SB_SB4_U134 ( .A1(R2_SB_SB4_n853), .A2(R2_SB_SB4_n829), .B1(
        R2_SB_SB4_n608), .B2(R2_SB_SB4_n826), .C1(R2_SB_SB4_n870), .C2(
        R2_SB_SB4_n831), .ZN(R2_SB_SB4_n465) );
  NOR3_X1 R2_SB_SB4_U133 ( .A1(R2_SB_SB4_n877), .A2(R2_SB_SB4_n638), .A3(
        R2_SB_SB4_n679), .ZN(R2_SB_SB4_n466) );
  INV_X1 R2_SB_SB4_U132 ( .A(R2_SB_SB4_n465), .ZN(R2_SB_SB4_n871) );
  OAI222_X1 R2_SB_SB4_U131 ( .A1(R2_SB_SB4_n871), .A2(R2_SB_SB4_n883), .B1(
        R2_SB_SB4_n849), .B2(R2_SB_SB4_n769), .C1(R2_SB_SB4_n466), .C2(
        R2_SB_SB4_n834), .ZN(R2_SB_SB4_n484) );
  INV_X1 R2_SB_SB4_U130 ( .A(R2_SB_SB4_n782), .ZN(R2_SB_SB4_n849) );
  NOR2_X1 R2_SB_SB4_U129 ( .A1(R2_SB_SB4_n830), .A2(R2_SB_SB4_n854), .ZN(
        R2_SB_SB4_n627) );
  NOR2_X1 R2_SB_SB4_U128 ( .A1(R2_SB_SB4_n881), .A2(R2_SB_SB4_n872), .ZN(
        R2_SB_SB4_n669) );
  INV_X1 R2_SB_SB4_U127 ( .A(R2_SB_SB4_n702), .ZN(R2_SB_SB4_n905) );
  NOR2_X1 R2_SB_SB4_U126 ( .A1(R2_SB_SB4_n453), .A2(R2_SB_SB4_n830), .ZN(
        R2_SB_SB4_n766) );
  NOR3_X1 R2_SB_SB4_U125 ( .A1(R2_SB_SB4_n828), .A2(R2_SB_SB4_n854), .A3(
        R2_SB_SB4_n908), .ZN(R2_SB_SB4_n673) );
  NOR2_X1 R2_SB_SB4_U124 ( .A1(R2_SB_SB4_n89), .A2(R2_SB_SB4_n830), .ZN(
        R2_SB_SB4_n771) );
  NOR2_X1 R2_SB_SB4_U123 ( .A1(R2_SB_SB4_n863), .A2(R2_SB_SB4_n843), .ZN(
        R2_SB_SB4_n778) );
  NOR2_X1 R2_SB_SB4_U122 ( .A1(R2_SB_SB4_n830), .A2(R2_SB_n290), .ZN(
        R2_SB_SB4_n779) );
  AOI21_X1 R2_SB_SB4_U121 ( .B1(R2_SB_SB4_n826), .B2(R2_SB_SB4_n833), .A(
        R2_SB_SB4_n800), .ZN(R2_SB_SB4_n549) );
  INV_X1 R2_SB_SB4_U120 ( .A(R2_SB_SB4_n549), .ZN(R2_SB_SB4_n902) );
  AND3_X1 R2_SB_SB4_U119 ( .A1(R2_SB_SB4_n548), .A2(R2_SB_SB4_n838), .A3(
        R2_SB_SB4_n849), .ZN(R2_SB_SB4_n550) );
  OR3_X1 R2_SB_SB4_U118 ( .A1(R2_SB_SB4_n864), .A2(R2_SB_SB4_n814), .A3(
        R2_SB_SB4_n890), .ZN(R2_SB_SB4_n815) );
  INV_X1 R2_SB_SB4_U117 ( .A(R2_SB_SB4_n519), .ZN(R2_SB_SB4_n886) );
  INV_X1 R2_SB_SB4_U116 ( .A(R2_SB_SB4_n790), .ZN(R2_SB_SB4_n866) );
  NAND2_X1 R2_SB_SB4_U115 ( .A1(R2_SB_SB4_n874), .A2(R2_SB_SB4_n901), .ZN(
        R2_SB_SB4_n728) );
  NAND2_X1 R2_SB_SB4_U114 ( .A1(R2_SB_SB4_n890), .A2(R2_SB_SB4_n874), .ZN(
        R2_SB_SB4_n536) );
  NAND2_X1 R2_SB_SB4_U113 ( .A1(R2_SB_SB4_n836), .A2(R2_SB_SB4_n826), .ZN(
        R2_SB_SB4_n723) );
  NAND2_X1 R2_SB_SB4_U112 ( .A1(R2_SB_SB4_n905), .A2(R2_SB_SB4_n875), .ZN(
        R2_SB_SB4_n589) );
  INV_X1 R2_SB_SB4_U111 ( .A(R2_SB_SB4_n627), .ZN(R2_SB_SB4_n856) );
  NAND2_X1 R2_SB_SB4_U110 ( .A1(R2_SB_SB4_n836), .A2(R2_SB_SB4_n829), .ZN(
        R2_SB_SB4_n748) );
  AND2_X1 R2_SB_SB4_U109 ( .A1(R2_SB_SB4_n766), .A2(R2_SB_SB4_n671), .ZN(
        R2_SB_SB4_n555) );
  INV_X1 R2_SB_SB4_U108 ( .A(R2_SB_SB4_n812), .ZN(R2_SB_SB4_n875) );
  OAI21_X1 R2_SB_SB4_U107 ( .B1(R2_SB_SB4_n847), .B2(R2_SB_SB4_n895), .A(
        R2_SB_SB4_n800), .ZN(R2_SB_SB4_n806) );
  NAND2_X1 R2_SB_SB4_U106 ( .A1(R2_SB_SB4_n628), .A2(R2_SB_SB4_n634), .ZN(
        R2_SB_SB4_n769) );
  NAND2_X1 R2_SB_SB4_U105 ( .A1(R2_SB_SB4_n507), .A2(R2_SB_SB4_n669), .ZN(
        R2_SB_SB4_n588) );
  INV_X1 R2_SB_SB4_U104 ( .A(R2_SB_SB4_n634), .ZN(R2_SB_SB4_n903) );
  INV_X1 R2_SB_SB4_U103 ( .A(R2_SB_SB4_n778), .ZN(R2_SB_SB4_n865) );
  NOR2_X1 R2_SB_SB4_U102 ( .A1(R2_SB_SB4_n730), .A2(R2_SB_SB4_n758), .ZN(
        R2_SB_SB4_n685) );
  AOI21_X1 R2_SB_SB4_U101 ( .B1(R2_SB_SB4_n588), .B2(R2_SB_SB4_n773), .A(
        R2_SB_SB4_n836), .ZN(R2_SB_SB4_n460) );
  AOI21_X1 R2_SB_SB4_U100 ( .B1(R2_SB_SB4_n802), .B2(R2_SB_SB4_n801), .A(
        R2_SB_SB4_n835), .ZN(R2_SB_SB4_n803) );
  INV_X1 R2_SB_SB4_U99 ( .A(R2_SB_SB4_n672), .ZN(R2_SB_SB4_n888) );
  NOR4_X1 R2_SB_SB4_U98 ( .A1(R2_SB_SB4_n675), .A2(R2_SB_SB4_n888), .A3(
        R2_SB_SB4_n674), .A4(R2_SB_SB4_n673), .ZN(R2_SB_SB4_n676) );
  NAND2_X1 R2_SB_SB4_U97 ( .A1(R2_SB_SB4_n778), .A2(R2_SB_SB4_n669), .ZN(
        R2_SB_SB4_n573) );
  INV_X1 R2_SB_SB4_U96 ( .A(R2_SB_SB4_n648), .ZN(R2_SB_SB4_n882) );
  NOR2_X1 R2_SB_SB4_U95 ( .A1(R2_SB_SB4_n849), .A2(R2_SB_SB4_n89), .ZN(
        R2_SB_SB4_n502) );
  NOR2_X1 R2_SB_SB4_U94 ( .A1(R2_SB_SB4_n851), .A2(R2_SB_n290), .ZN(
        R2_SB_SB4_n470) );
  NOR2_X1 R2_SB_SB4_U93 ( .A1(R2_SB_SB4_n853), .A2(R2_SB_SB4_n903), .ZN(
        R2_SB_SB4_n514) );
  INV_X1 R2_SB_SB4_U92 ( .A(R2_SB_SB4_n604), .ZN(R2_SB_SB4_n844) );
  NOR2_X1 R2_SB_SB4_U91 ( .A1(R2_SB_SB4_n862), .A2(R2_SB_SB4_n883), .ZN(
        R2_SB_SB4_n534) );
  INV_X1 R2_SB_SB4_U90 ( .A(R2_SB_SB4_n603), .ZN(R2_SB_SB4_n848) );
  INV_X1 R2_SB_SB4_U89 ( .A(R2_SB_SB4_n802), .ZN(R2_SB_SB4_n877) );
  NOR2_X1 R2_SB_SB4_U88 ( .A1(R2_SB_SB4_n905), .A2(R2_SB_SB4_n866), .ZN(
        R2_SB_SB4_n671) );
  OAI22_X1 R2_SB_SB4_U87 ( .A1(R2_SB_SB4_n730), .A2(R2_SB_SB4_n905), .B1(
        R2_SB_SB4_n901), .B2(R2_SB_SB4_n851), .ZN(R2_SB_SB4_n462) );
  OAI22_X1 R2_SB_SB4_U86 ( .A1(R2_SB_SB4_n875), .A2(R2_SB_SB4_n833), .B1(
        R2_SB_SB4_n874), .B2(R2_SB_SB4_n832), .ZN(R2_SB_SB4_n804) );
  OAI22_X1 R2_SB_SB4_U85 ( .A1(R2_SB_SB4_n665), .A2(R2_SB_SB4_n892), .B1(
        R2_SB_SB4_n841), .B2(R2_SB_SB4_n801), .ZN(R2_SB_SB4_n666) );
  INV_X1 R2_SB_SB4_U84 ( .A(R2_SB_SB4_n758), .ZN(R2_SB_SB4_n847) );
  AOI21_X1 R2_SB_SB4_U83 ( .B1(R2_SB_SB4_n868), .B2(R2_SB_SB4_n845), .A(
        R2_SB_SB4_n785), .ZN(R2_SB_SB4_n687) );
  OAI22_X1 R2_SB_SB4_U82 ( .A1(R2_SB_SB4_n831), .A2(R2_SB_SB4_n895), .B1(
        R2_SB_n289), .B2(R2_SB_SB4_n648), .ZN(R2_SB_SB4_n532) );
  AOI22_X1 R2_SB_SB4_U81 ( .A1(R2_SB_SB4_n758), .A2(R2_SB_n290), .B1(
        R2_SB_SB4_n771), .B2(R2_SB_SB4_n452), .ZN(R2_SB_SB4_n699) );
  INV_X1 R2_SB_SB4_U80 ( .A(R2_SB_SB4_n771), .ZN(R2_SB_SB4_n831) );
  NOR2_X1 R2_SB_SB4_U79 ( .A1(R2_SB_SB4_n842), .A2(R2_SB_SB4_n898), .ZN(
        R2_SB_SB4_n675) );
  NOR2_X1 R2_SB_SB4_U78 ( .A1(R2_SB_SB4_n868), .A2(R2_SB_SB4_n890), .ZN(
        R2_SB_SB4_n576) );
  NOR2_X1 R2_SB_SB4_U77 ( .A1(R2_SB_SB4_n774), .A2(R2_SB_SB4_n890), .ZN(
        R2_SB_SB4_n565) );
  NOR2_X1 R2_SB_SB4_U76 ( .A1(R2_SB_SB4_n845), .A2(R2_SB_SB4_n89), .ZN(
        R2_SB_SB4_n725) );
  NOR2_X1 R2_SB_SB4_U75 ( .A1(R2_SB_SB4_n853), .A2(R2_SB_SB4_n890), .ZN(
        R2_SB_SB4_n633) );
  NOR2_X1 R2_SB_SB4_U74 ( .A1(R2_SB_SB4_n868), .A2(R2_SB_SB4_n905), .ZN(
        R2_SB_SB4_n754) );
  NOR2_X1 R2_SB_SB4_U73 ( .A1(R2_SB_SB4_n869), .A2(R2_SB_SB4_n905), .ZN(
        R2_SB_SB4_n698) );
  NOR2_X1 R2_SB_SB4_U72 ( .A1(R2_SB_SB4_n898), .A2(R2_SB_SB4_n845), .ZN(
        R2_SB_SB4_n756) );
  NOR2_X1 R2_SB_SB4_U71 ( .A1(R2_SB_SB4_n774), .A2(R2_SB_SB4_n905), .ZN(
        R2_SB_SB4_n638) );
  NOR2_X1 R2_SB_SB4_U70 ( .A1(R2_SB_SB4_n870), .A2(R2_SB_SB4_n890), .ZN(
        R2_SB_SB4_n727) );
  OAI22_X1 R2_SB_SB4_U69 ( .A1(R2_SB_SB4_n453), .A2(R2_SB_SB4_n879), .B1(
        R2_SB_SB4_n89), .B2(R2_SB_SB4_n880), .ZN(R2_SB_SB4_n538) );
  AOI211_X1 R2_SB_SB4_U68 ( .C1(R2_SB_SB4_n576), .C2(R2_SB_SB4_n89), .A(
        R2_SB_SB4_n538), .B(R2_SB_SB4_n722), .ZN(R2_SB_SB4_n543) );
  INV_X1 R2_SB_SB4_U67 ( .A(R2_SB_SB4_n779), .ZN(R2_SB_SB4_n833) );
  NOR3_X1 R2_SB_SB4_U66 ( .A1(R2_SB_SB4_n841), .A2(R2_SB_SB4_n858), .A3(
        R2_SB_SB4_n874), .ZN(R2_SB_SB4_n521) );
  INV_X1 R2_SB_SB4_U65 ( .A(R2_SB_SB4_n766), .ZN(R2_SB_SB4_n835) );
  NOR2_X1 R2_SB_SB4_U64 ( .A1(R2_SB_SB4_n838), .A2(R2_SB_SB4_n453), .ZN(
        R2_SB_SB4_n742) );
  INV_X1 R2_SB_SB4_U63 ( .A(R2_SB_SB4_n730), .ZN(R2_SB_SB4_n858) );
  NOR2_X1 R2_SB_SB4_U62 ( .A1(R2_SB_SB4_n878), .A2(R2_SB_SB4_n869), .ZN(
        R2_SB_SB4_n713) );
  NOR2_X1 R2_SB_SB4_U61 ( .A1(R2_SB_SB4_n833), .A2(R2_SB_SB4_n453), .ZN(
        R2_SB_SB4_n799) );
  AOI22_X1 R2_SB_SB4_U60 ( .A1(R2_SB_SB4_n877), .A2(R2_SB_SB4_n452), .B1(
        R2_SB_SB4_n781), .B2(R2_SB_SB4_n669), .ZN(R2_SB_SB4_n500) );
  OAI211_X1 R2_SB_SB4_U59 ( .C1(R2_SB_SB4_n89), .C2(R2_SB_SB4_n893), .A(
        R2_SB_SB4_n907), .B(R2_SB_SB4_n500), .ZN(R2_SB_SB4_n501) );
  AOI222_X1 R2_SB_SB4_U58 ( .A1(R2_SB_SB4_n591), .A2(R2_SB_SB4_n748), .B1(
        R2_SB_SB4_n502), .B2(R2_SB_SB4_n679), .C1(R2_SB_SB4_n758), .C2(
        R2_SB_SB4_n501), .ZN(R2_SB_SB4_n526) );
  OAI222_X1 R2_SB_SB4_U57 ( .A1(R2_SB_SB4_n845), .A2(R2_SB_SB4_n880), .B1(
        R2_SB_SB4_n835), .B2(R2_SB_SB4_n898), .C1(R2_SB_SB4_n836), .C2(
        R2_SB_SB4_n894), .ZN(R2_SB_SB4_n602) );
  NOR2_X1 R2_SB_SB4_U56 ( .A1(R2_SB_SB4_n883), .A2(R2_SB_SB4_n869), .ZN(
        R2_SB_SB4_n755) );
  NOR2_X1 R2_SB_SB4_U55 ( .A1(R2_SB_SB4_n862), .A2(R2_SB_SB4_n890), .ZN(
        R2_SB_SB4_n753) );
  NOR2_X1 R2_SB_SB4_U54 ( .A1(R2_SB_SB4_n862), .A2(R2_SB_SB4_n905), .ZN(
        R2_SB_SB4_n759) );
  NOR2_X1 R2_SB_SB4_U53 ( .A1(R2_SB_SB4_n862), .A2(R2_SB_SB4_n878), .ZN(
        R2_SB_SB4_n591) );
  NOR2_X1 R2_SB_SB4_U52 ( .A1(R2_SB_SB4_n869), .A2(R2_SB_SB4_n890), .ZN(
        R2_SB_SB4_n679) );
  INV_X1 R2_SB_SB4_U51 ( .A(R2_SB_SB4_n669), .ZN(R2_SB_SB4_n890) );
  NOR2_X2 R2_SB_SB4_U50 ( .A1(R2_SB_SB4_n89), .A2(R2_SB_SB4_n453), .ZN(
        R2_SB_SB4_n781) );
  NOR2_X2 R2_SB_SB4_U49 ( .A1(R2_SB_SB4_n89), .A2(R2_SB_SB4_n452), .ZN(
        R2_SB_SB4_n684) );
  NOR3_X1 R2_SB_SB4_U48 ( .A1(R2_SB_SB4_n878), .A2(R2_SB_SB4_n866), .A3(
        R2_SB_SB4_n838), .ZN(R2_SB_SB4_n674) );
  NOR2_X1 R2_SB_SB4_U47 ( .A1(R2_SB_SB4_n840), .A2(R2_SB_SB4_n452), .ZN(
        R2_SB_SB4_n747) );
  NOR2_X1 R2_SB_SB4_U46 ( .A1(R2_SB_SB4_n453), .A2(R2_SB_n290), .ZN(
        R2_SB_SB4_n810) );
  INV_X1 R2_SB_SB4_U45 ( .A(R2_SB_SB4_n633), .ZN(R2_SB_SB4_n891) );
  INV_X1 R2_SB_SB4_U44 ( .A(R2_SB_SB4_n534), .ZN(R2_SB_SB4_n885) );
  INV_X1 R2_SB_SB4_U43 ( .A(R2_SB_SB4_n470), .ZN(R2_SB_SB4_n852) );
  INV_X1 R2_SB_SB4_U42 ( .A(R2_SB_SB4_n502), .ZN(R2_SB_SB4_n850) );
  INV_X1 R2_SB_SB4_U41 ( .A(R2_SB_SB4_n514), .ZN(R2_SB_SB4_n904) );
  INV_X1 R2_SB_SB4_U40 ( .A(R2_SB_SB4_n698), .ZN(R2_SB_SB4_n906) );
  INV_X1 R2_SB_SB4_U39 ( .A(R2_SB_SB4_n638), .ZN(R2_SB_SB4_n908) );
  INV_X1 R2_SB_SB4_U38 ( .A(R2_SB_SB4_n565), .ZN(R2_SB_SB4_n892) );
  INV_X1 R2_SB_SB4_U37 ( .A(R2_SB_SB4_n753), .ZN(R2_SB_SB4_n893) );
  INV_X1 R2_SB_SB4_U36 ( .A(R2_SB_SB4_n727), .ZN(R2_SB_SB4_n894) );
  INV_X1 R2_SB_SB4_U35 ( .A(R2_SB_SB4_n755), .ZN(R2_SB_SB4_n884) );
  INV_X1 R2_SB_SB4_U34 ( .A(R2_SB_SB4_n799), .ZN(R2_SB_SB4_n834) );
  NAND2_X1 R2_SB_SB4_U33 ( .A1(R2_SB_SB4_n781), .A2(R2_SB_SB4_n671), .ZN(
        R2_SB_SB4_n716) );
  INV_X1 R2_SB_SB4_U32 ( .A(R2_SB_SB4_n588), .ZN(R2_SB_SB4_n900) );
  INV_X1 R2_SB_SB4_U31 ( .A(R2_SB_SB4_n759), .ZN(R2_SB_SB4_n907) );
  INV_X1 R2_SB_SB4_U30 ( .A(R2_SB_SB4_n747), .ZN(R2_SB_SB4_n841) );
  INV_X1 R2_SB_SB4_U29 ( .A(R2_SB_SB4_n713), .ZN(R2_SB_SB4_n879) );
  INV_X1 R2_SB_SB4_U28 ( .A(R2_SB_SB4_n591), .ZN(R2_SB_SB4_n880) );
  INV_X1 R2_SB_SB4_U27 ( .A(R2_SB_SB4_n742), .ZN(R2_SB_SB4_n839) );
  AOI21_X1 R2_SB_SB4_U26 ( .B1(R2_SB_SB4_n848), .B2(R2_SB_SB4_n852), .A(
        R2_SB_SB4_n910), .ZN(R2_SB_SB4_n461) );
  AOI21_X1 R2_SB_SB4_U25 ( .B1(R2_SB_SB4_n831), .B2(R2_SB_SB4_n835), .A(
        R2_SB_SB4_n890), .ZN(R2_SB_SB4_n796) );
  INV_X1 R2_SB_SB4_U24 ( .A(R2_SB_SB4_n684), .ZN(R2_SB_SB4_n827) );
  AOI22_X1 R2_SB_SB4_U23 ( .A1(R2_SB_SB4_n877), .A2(R2_SB_n290), .B1(
        R2_SB_SB4_n713), .B2(R2_SB_SB4_n828), .ZN(R2_SB_SB4_n649) );
  INV_X1 R2_SB_SB4_U22 ( .A(R2_SB_SB4_n754), .ZN(R2_SB_SB4_n910) );
  INV_X1 R2_SB_SB4_U21 ( .A(R2_SB_SB4_n781), .ZN(R2_SB_SB4_n828) );
  INV_X1 R2_SB_SB4_U20 ( .A(R2_SB_SB4_n576), .ZN(R2_SB_SB4_n898) );
  INV_X1 R2_SB_SB4_U19 ( .A(R2_SB_SB4_n679), .ZN(R2_SB_SB4_n895) );
  NOR2_X1 R2_SB_SB4_U18 ( .A1(R2_SB_SB4_n831), .A2(R2_SB_SB4_n452), .ZN(
        R2_SB_SB4_n708) );
  OAI221_X1 R2_SB_SB4_U17 ( .B1(R2_SB_n290), .B2(R2_SB_SB4_n906), .C1(
        R2_SB_SB4_n890), .C2(R2_SB_SB4_n826), .A(R2_SB_SB4_n769), .ZN(
        R2_SB_SB4_n590) );
  NOR2_X1 R2_SB_SB4_U16 ( .A1(R2_SB_SB4_n895), .A2(R2_SB_SB4_n452), .ZN(
        R2_SB_SB4_n722) );
  INV_X1 R2_SB_SB4_U15 ( .A(R2_SB_SB4_n810), .ZN(R2_SB_SB4_n829) );
  NOR2_X1 R2_SB_SB4_U14 ( .A1(R2_SB_n289), .A2(R2_SB_n290), .ZN(R2_SB_SB4_n628) );
  INV_X1 R2_SB_SB4_U13 ( .A(R2_SB_SB4_n708), .ZN(R2_SB_SB4_n832) );
  INV_X1 R2_SB_SB4_U12 ( .A(R2_SB_SB4_n628), .ZN(R2_SB_SB4_n826) );
  NOR2_X1 R2_SB_SB4_U11 ( .A1(R2_SB_SB4_n863), .A2(R2_SB_n293), .ZN(
        R2_SB_SB4_n744) );
  NOR2_X1 R2_SB_SB4_U10 ( .A1(R2_SB_SB4_n881), .A2(R2_SB_n295), .ZN(
        R2_SB_SB4_n772) );
  NOR2_X1 R2_SB_SB4_U9 ( .A1(R2_SB_SB4_n89), .A2(R2_SB_n291), .ZN(
        R2_SB_SB4_n791) );
  NOR2_X1 R2_SB_SB4_U8 ( .A1(R2_SB_SB4_n872), .A2(R2_SB_n296), .ZN(
        R2_SB_SB4_n752) );
  NOR2_X1 R2_SB_SB4_U7 ( .A1(R2_SB_SB4_n854), .A2(R2_SB_SB4_n843), .ZN(
        R2_SB_SB4_n730) );
  NOR2_X1 R2_SB_SB4_U6 ( .A1(R2_SB_SB4_n843), .A2(R2_SB_n294), .ZN(
        R2_SB_SB4_n780) );
  NOR2_X1 R2_SB_SB4_U5 ( .A1(R2_SB_n291), .A2(R2_SB_n292), .ZN(R2_SB_SB4_n743)
         );
  INV_X1 R2_SB_SB4_U4 ( .A(R2_SB_n292), .ZN(R2_SB_SB4_n843) );
  NOR2_X1 R2_SB_SB4_U3 ( .A1(R2_SB_SB4_n453), .A2(R2_SB_n291), .ZN(
        R2_SB_SB4_n696) );
  NOR2_X1 R2_SB_SB4_U2 ( .A1(R2_SB_SB4_n881), .A2(R2_SB_n294), .ZN(
        R2_SB_SB4_n798) );
  NOR2_X1 R2_SB_SB4_U1 ( .A1(R2_SB_SB4_n843), .A2(R2_SB_n293), .ZN(
        R2_SB_SB4_n789) );
  NAND3_X1 R2_SB_SB4_U464 ( .A1(R2_SB_SB4_n772), .A2(R2_SB_SB4_n670), .A3(
        R2_SB_SB4_n794), .ZN(R2_SB_SB4_n519) );
  OAI33_X1 R2_SB_SB4_U463 ( .A1(R2_SB_SB4_n838), .A2(R2_SB_SB4_n858), .A3(
        R2_SB_SB4_n905), .B1(R2_SB_SB4_n853), .B2(R2_SB_SB4_n830), .B3(
        R2_SB_SB4_n874), .ZN(R2_SB_SB4_n467) );
  NAND3_X1 R2_SB_SB4_U462 ( .A1(R2_SB_SB4_n507), .A2(R2_SB_SB4_n702), .A3(
        R2_SB_SB4_n758), .ZN(R2_SB_SB4_n677) );
  OAI33_X1 R2_SB_SB4_U461 ( .A1(R2_SB_SB4_n828), .A2(R2_SB_n296), .A3(
        R2_SB_n291), .B1(R2_SB_SB4_n472), .B2(R2_SB_SB4_n854), .B3(
        R2_SB_SB4_n829), .ZN(R2_SB_SB4_n473) );
  NAND4_X1 R2_SB_SB4_U460 ( .A1(R2_SB_SB4_n488), .A2(R2_SB_SB4_n487), .A3(
        R2_SB_SB4_n486), .A4(R2_SB_SB4_n485), .ZN(R2_SB_n[281]) );
  NAND3_X1 R2_SB_SB4_U459 ( .A1(R2_SB_SB4_n781), .A2(R2_SB_n291), .A3(
        R2_SB_SB4_n798), .ZN(R2_SB_SB4_n494) );
  NAND4_X1 R2_SB_SB4_U458 ( .A1(R2_SB_SB4_n743), .A2(R2_SB_SB4_n628), .A3(
        R2_SB_SB4_n767), .A4(R2_SB_n296), .ZN(R2_SB_SB4_n493) );
  NAND3_X1 R2_SB_SB4_U457 ( .A1(R2_SB_SB4_n813), .A2(R2_SB_SB4_n830), .A3(
        R2_SB_SB4_n684), .ZN(R2_SB_SB4_n492) );
  NAND3_X1 R2_SB_SB4_U456 ( .A1(R2_SB_SB4_n494), .A2(R2_SB_SB4_n493), .A3(
        R2_SB_SB4_n492), .ZN(R2_SB_SB4_n498) );
  NAND3_X1 R2_SB_SB4_U455 ( .A1(R2_SB_SB4_n844), .A2(R2_SB_SB4_n836), .A3(
        R2_SB_SB4_n548), .ZN(R2_SB_SB4_n506) );
  OAI33_X1 R2_SB_SB4_U454 ( .A1(R2_SB_SB4_n827), .A2(R2_SB_SB4_n856), .A3(
        R2_SB_SB4_n903), .B1(R2_SB_SB4_n898), .B2(R2_SB_SB4_n843), .B3(
        R2_SB_SB4_n826), .ZN(R2_SB_SB4_n515) );
  NAND3_X1 R2_SB_SB4_U453 ( .A1(R2_SB_SB4_n671), .A2(R2_SB_SB4_n453), .A3(
        R2_SB_n291), .ZN(R2_SB_SB4_n816) );
  NAND3_X1 R2_SB_SB4_U452 ( .A1(R2_SB_SB4_n670), .A2(R2_SB_SB4_n669), .A3(
        R2_SB_SB4_n779), .ZN(R2_SB_SB4_n672) );
  NAND3_X1 R2_SB_SB4_U451 ( .A1(R2_SB_SB4_n816), .A2(R2_SB_SB4_n519), .A3(
        R2_SB_SB4_n672), .ZN(R2_SB_SB4_n522) );
  OAI33_X1 R2_SB_SB4_U450 ( .A1(R2_SB_SB4_n832), .A2(R2_SB_SB4_n864), .A3(
        R2_SB_SB4_n890), .B1(R2_SB_SB4_n829), .B2(R2_SB_n296), .B3(
        R2_SB_SB4_n866), .ZN(R2_SB_SB4_n520) );
  NAND4_X1 R2_SB_SB4_U449 ( .A1(R2_SB_SB4_n527), .A2(R2_SB_SB4_n526), .A3(
        R2_SB_SB4_n525), .A4(R2_SB_SB4_n524), .ZN(R2_SB_n[282]) );
  NAND3_X1 R2_SB_SB4_U448 ( .A1(R2_SB_SB4_n744), .A2(R2_SB_SB4_n603), .A3(
        R2_SB_SB4_n696), .ZN(R2_SB_SB4_n546) );
  NAND3_X1 R2_SB_SB4_U447 ( .A1(R2_SB_SB4_n684), .A2(R2_SB_SB4_n854), .A3(
        R2_SB_SB4_n709), .ZN(R2_SB_SB4_n582) );
  OAI33_X1 R2_SB_SB4_U446 ( .A1(R2_SB_SB4_n859), .A2(R2_SB_SB4_n830), .A3(
        R2_SB_SB4_n901), .B1(R2_SB_SB4_n876), .B2(R2_SB_n290), .B3(
        R2_SB_SB4_n685), .ZN(R2_SB_SB4_n557) );
  NAND4_X1 R2_SB_SB4_U445 ( .A1(R2_SB_SB4_n561), .A2(R2_SB_SB4_n560), .A3(
        R2_SB_SB4_n559), .A4(R2_SB_SB4_n558), .ZN(R2_SB_n[283]) );
  NAND3_X1 R2_SB_SB4_U444 ( .A1(R2_SB_SB4_n830), .A2(R2_SB_SB4_n872), .A3(
        R2_SB_SB4_n709), .ZN(R2_SB_SB4_n566) );
  NAND4_X1 R2_SB_SB4_U443 ( .A1(R2_SB_SB4_n566), .A2(R2_SB_SB4_n894), .A3(
        R2_SB_SB4_n800), .A4(R2_SB_SB4_n648), .ZN(R2_SB_SB4_n569) );
  NAND3_X1 R2_SB_SB4_U442 ( .A1(R2_SB_n289), .A2(R2_SB_n292), .A3(
        R2_SB_SB4_n744), .ZN(R2_SB_SB4_n659) );
  NAND3_X1 R2_SB_SB4_U441 ( .A1(R2_SB_SB4_n758), .A2(R2_SB_SB4_n854), .A3(
        R2_SB_SB4_n709), .ZN(R2_SB_SB4_n587) );
  NAND3_X1 R2_SB_SB4_U440 ( .A1(R2_SB_SB4_n743), .A2(R2_SB_n289), .A3(
        R2_SB_SB4_n882), .ZN(R2_SB_SB4_n592) );
  NAND4_X1 R2_SB_SB4_U439 ( .A1(R2_SB_SB4_n601), .A2(R2_SB_SB4_n600), .A3(
        R2_SB_SB4_n599), .A4(R2_SB_SB4_n598), .ZN(R2_SB_n[284]) );
  NAND4_X1 R2_SB_SB4_U438 ( .A1(R2_SB_SB4_n645), .A2(R2_SB_SB4_n644), .A3(
        R2_SB_SB4_n643), .A4(R2_SB_SB4_n642), .ZN(R2_SB_n[285]) );
  NAND3_X1 R2_SB_SB4_U437 ( .A1(R2_SB_SB4_n684), .A2(R2_SB_SB4_n843), .A3(
        R2_SB_SB4_n744), .ZN(R2_SB_SB4_n660) );
  NAND3_X1 R2_SB_SB4_U436 ( .A1(R2_SB_n289), .A2(R2_SB_SB4_n854), .A3(
        R2_SB_SB4_n792), .ZN(R2_SB_SB4_n658) );
  NAND4_X1 R2_SB_SB4_U435 ( .A1(R2_SB_SB4_n660), .A2(R2_SB_SB4_n659), .A3(
        R2_SB_SB4_n658), .A4(R2_SB_SB4_n657), .ZN(R2_SB_SB4_n668) );
  OAI33_X1 R2_SB_SB4_U434 ( .A1(R2_SB_SB4_n862), .A2(R2_SB_n296), .A3(
        R2_SB_SB4_n847), .B1(R2_SB_SB4_n903), .B2(R2_SB_SB4_n858), .B3(
        R2_SB_SB4_n830), .ZN(R2_SB_SB4_n661) );
  NAND3_X1 R2_SB_SB4_U433 ( .A1(R2_SB_SB4_n670), .A2(R2_SB_SB4_n669), .A3(
        R2_SB_SB4_n766), .ZN(R2_SB_SB4_n717) );
  NAND4_X1 R2_SB_SB4_U432 ( .A1(R2_SB_SB4_n717), .A2(R2_SB_SB4_n716), .A3(
        R2_SB_SB4_n677), .A4(R2_SB_SB4_n676), .ZN(R2_SB_SB4_n689) );
  OAI33_X1 R2_SB_SB4_U431 ( .A1(R2_SB_SB4_n839), .A2(R2_SB_SB4_n870), .A3(
        R2_SB_SB4_n883), .B1(R2_SB_SB4_n827), .B2(R2_SB_SB4_n685), .B3(
        R2_SB_SB4_n903), .ZN(R2_SB_SB4_n686) );
  NAND4_X1 R2_SB_SB4_U430 ( .A1(R2_SB_SB4_n693), .A2(R2_SB_SB4_n692), .A3(
        R2_SB_SB4_n691), .A4(R2_SB_SB4_n690), .ZN(R2_SB_n[286]) );
  NAND3_X1 R2_SB_SB4_U429 ( .A1(R2_SB_SB4_n845), .A2(R2_SB_SB4_n838), .A3(
        R2_SB_SB4_n829), .ZN(R2_SB_SB4_n703) );
  OAI33_X1 R2_SB_SB4_U428 ( .A1(R2_SB_SB4_n876), .A2(R2_SB_n289), .A3(
        R2_SB_SB4_n830), .B1(R2_SB_SB4_n705), .B2(R2_SB_SB4_n835), .B3(
        R2_SB_SB4_n901), .ZN(R2_SB_SB4_n706) );
  NAND3_X1 R2_SB_SB4_U427 ( .A1(R2_SB_n293), .A2(R2_SB_SB4_n714), .A3(
        R2_SB_n296), .ZN(R2_SB_SB4_n715) );
  NAND3_X1 R2_SB_SB4_U426 ( .A1(R2_SB_SB4_n717), .A2(R2_SB_SB4_n716), .A3(
        R2_SB_SB4_n715), .ZN(R2_SB_SB4_n737) );
  NAND4_X1 R2_SB_SB4_U425 ( .A1(R2_SB_SB4_n741), .A2(R2_SB_SB4_n740), .A3(
        R2_SB_SB4_n739), .A4(R2_SB_SB4_n738), .ZN(R2_SB_n[287]) );
  NAND3_X1 R2_SB_SB4_U424 ( .A1(R2_SB_n296), .A2(R2_SB_SB4_n854), .A3(
        R2_SB_SB4_n795), .ZN(R2_SB_SB4_n762) );
  NAND3_X1 R2_SB_SB4_U423 ( .A1(R2_SB_SB4_n763), .A2(R2_SB_SB4_n762), .A3(
        R2_SB_SB4_n761), .ZN(R2_SB_SB4_n764) );
  NAND3_X1 R2_SB_SB4_U422 ( .A1(R2_SB_n295), .A2(R2_SB_SB4_n854), .A3(
        R2_SB_SB4_n771), .ZN(R2_SB_SB4_n777) );
  NAND3_X1 R2_SB_SB4_U421 ( .A1(R2_SB_SB4_n817), .A2(R2_SB_SB4_n816), .A3(
        R2_SB_SB4_n815), .ZN(R2_SB_SB4_n820) );
  NAND4_X1 R2_SB_SB4_U420 ( .A1(R2_SB_SB4_n825), .A2(R2_SB_SB4_n824), .A3(
        R2_SB_SB4_n823), .A4(R2_SB_SB4_n822), .ZN(R2_SB_n[288]) );
  NOR2_X2 R2_SB_SB4_U264 ( .A1(R2_SB_SB4_n830), .A2(R2_SB_SB4_n843), .ZN(
        R2_SB_SB4_n758) );
  BUF_X1 R2_SR_U128 ( .A(R2_n1472), .Z(R2_n1280) );
  BUF_X1 R2_SR_U127 ( .A(R2_n1471), .Z(R2_n1279) );
  BUF_X1 R2_SR_U126 ( .A(R2_n1470), .Z(R2_n1278) );
  BUF_X1 R2_SR_U125 ( .A(R2_n1469), .Z(R2_n1277) );
  BUF_X1 R2_SR_U124 ( .A(R2_n1468), .Z(R2_n1276) );
  BUF_X1 R2_SR_U123 ( .A(R2_n1467), .Z(R2_n1275) );
  BUF_X1 R2_SR_U122 ( .A(R2_n1466), .Z(R2_n1274) );
  BUF_X1 R2_SR_U121 ( .A(R2_n1433), .Z(R2_n1273) );
  BUF_X1 R2_SR_U120 ( .A(R2_n1432), .Z(R2_n1272) );
  BUF_X1 R2_SR_U119 ( .A(R2_n1431), .Z(R2_n1271) );
  BUF_X1 R2_SR_U118 ( .A(R2_n1430), .Z(R2_n1270) );
  BUF_X1 R2_SR_U117 ( .A(R2_n1429), .Z(R2_n1269) );
  BUF_X1 R2_SR_U116 ( .A(R2_n1428), .Z(R2_n1268) );
  BUF_X1 R2_SR_U115 ( .A(R2_n1427), .Z(R2_n1267) );
  BUF_X1 R2_SR_U114 ( .A(R2_n1426), .Z(R2_n1266) );
  BUF_X1 R2_SR_U113 ( .A(R2_n1393), .Z(R2_n1265) );
  BUF_X1 R2_SR_U112 ( .A(R2_n1392), .Z(R2_n1264) );
  BUF_X1 R2_SR_U111 ( .A(R2_n1391), .Z(R2_n1263) );
  BUF_X1 R2_SR_U110 ( .A(R2_n1390), .Z(R2_n1262) );
  BUF_X1 R2_SR_U109 ( .A(R2_n1389), .Z(R2_n1261) );
  BUF_X1 R2_SR_U108 ( .A(R2_n1388), .Z(R2_n1260) );
  BUF_X1 R2_SR_U107 ( .A(R2_n1387), .Z(R2_n1259) );
  BUF_X1 R2_SR_U106 ( .A(R2_n1386), .Z(R2_n1258) );
  BUF_X1 R2_SR_U105 ( .A(R2_n1473), .Z(R2_n1281) );
  BUF_X1 R2_SR_U104 ( .A(R2_n1506), .Z(R2_n1282) );
  BUF_X1 R2_SR_U103 ( .A(R2_n1507), .Z(R2_n1283) );
  BUF_X1 R2_SR_U102 ( .A(R2_n1508), .Z(R2_n1284) );
  BUF_X1 R2_SR_U101 ( .A(R2_n1509), .Z(R2_n1285) );
  BUF_X1 R2_SR_U100 ( .A(R2_n1510), .Z(R2_n1286) );
  BUF_X1 R2_SR_U99 ( .A(R2_n1511), .Z(R2_n1287) );
  BUF_X1 R2_SR_U98 ( .A(R2_n1512), .Z(R2_n1288) );
  BUF_X1 R2_SR_U97 ( .A(R2_n1513), .Z(R2_n1289) );
  BUF_X1 R2_SR_U96 ( .A(R2_n1418), .Z(R2_n1290) );
  BUF_X1 R2_SR_U95 ( .A(R2_n1419), .Z(R2_n1291) );
  BUF_X1 R2_SR_U94 ( .A(R2_n1420), .Z(R2_n1292) );
  BUF_X1 R2_SR_U93 ( .A(R2_n1421), .Z(R2_n1293) );
  BUF_X1 R2_SR_U92 ( .A(R2_n1422), .Z(R2_n1294) );
  BUF_X1 R2_SR_U91 ( .A(R2_n1423), .Z(R2_n1295) );
  BUF_X1 R2_SR_U90 ( .A(R2_n1424), .Z(R2_n1296) );
  BUF_X1 R2_SR_U89 ( .A(R2_n1425), .Z(R2_n1297) );
  BUF_X1 R2_SR_U88 ( .A(R2_n1458), .Z(R2_n1298) );
  BUF_X1 R2_SR_U87 ( .A(R2_n1459), .Z(R2_n1299) );
  BUF_X1 R2_SR_U86 ( .A(R2_n1460), .Z(R2_n1300) );
  BUF_X1 R2_SR_U85 ( .A(R2_n1461), .Z(R2_n1301) );
  BUF_X1 R2_SR_U84 ( .A(R2_n1462), .Z(R2_n1302) );
  BUF_X1 R2_SR_U83 ( .A(R2_n1463), .Z(R2_n1303) );
  BUF_X1 R2_SR_U82 ( .A(R2_n1464), .Z(R2_n1304) );
  BUF_X1 R2_SR_U81 ( .A(R2_n1465), .Z(R2_n1305) );
  BUF_X1 R2_SR_U80 ( .A(R2_n1498), .Z(R2_n1306) );
  BUF_X1 R2_SR_U79 ( .A(R2_n1499), .Z(R2_n1307) );
  BUF_X1 R2_SR_U78 ( .A(R2_n1500), .Z(R2_n1308) );
  BUF_X1 R2_SR_U77 ( .A(R2_n1501), .Z(R2_n1309) );
  BUF_X1 R2_SR_U76 ( .A(R2_n1502), .Z(R2_n1310) );
  BUF_X1 R2_SR_U75 ( .A(R2_n1503), .Z(R2_n1311) );
  BUF_X1 R2_SR_U74 ( .A(R2_n1504), .Z(R2_n1312) );
  BUF_X1 R2_SR_U73 ( .A(R2_n1505), .Z(R2_n1313) );
  BUF_X1 R2_SR_U72 ( .A(R2_n1410), .Z(R2_n1314) );
  BUF_X1 R2_SR_U71 ( .A(R2_n1411), .Z(R2_n1315) );
  BUF_X1 R2_SR_U70 ( .A(R2_n1412), .Z(R2_n1316) );
  BUF_X1 R2_SR_U69 ( .A(R2_n1413), .Z(R2_n1317) );
  BUF_X1 R2_SR_U68 ( .A(R2_n1414), .Z(R2_n1318) );
  BUF_X1 R2_SR_U67 ( .A(R2_n1415), .Z(R2_n1319) );
  BUF_X1 R2_SR_U66 ( .A(R2_n1416), .Z(R2_n1320) );
  BUF_X1 R2_SR_U65 ( .A(R2_n1417), .Z(R2_n1321) );
  BUF_X1 R2_SR_U64 ( .A(R2_n1450), .Z(R2_n1322) );
  BUF_X1 R2_SR_U63 ( .A(R2_n1451), .Z(R2_n1323) );
  BUF_X1 R2_SR_U62 ( .A(R2_n1452), .Z(R2_n1324) );
  BUF_X1 R2_SR_U61 ( .A(R2_n1453), .Z(R2_n1325) );
  BUF_X1 R2_SR_U60 ( .A(R2_n1454), .Z(R2_n1326) );
  BUF_X1 R2_SR_U59 ( .A(R2_n1455), .Z(R2_n1327) );
  BUF_X1 R2_SR_U58 ( .A(R2_n1456), .Z(R2_n1328) );
  BUF_X1 R2_SR_U57 ( .A(R2_n1457), .Z(R2_n1329) );
  BUF_X1 R2_SR_U56 ( .A(R2_n1490), .Z(R2_n1330) );
  BUF_X1 R2_SR_U55 ( .A(R2_n1491), .Z(R2_n1331) );
  BUF_X1 R2_SR_U54 ( .A(R2_n1492), .Z(R2_n1332) );
  BUF_X1 R2_SR_U53 ( .A(R2_n1493), .Z(R2_n1333) );
  BUF_X1 R2_SR_U52 ( .A(R2_n1494), .Z(R2_n1334) );
  BUF_X1 R2_SR_U51 ( .A(R2_n1495), .Z(R2_n1335) );
  BUF_X1 R2_SR_U50 ( .A(R2_n1496), .Z(R2_n1336) );
  BUF_X1 R2_SR_U49 ( .A(R2_n1497), .Z(R2_n1337) );
  BUF_X1 R2_SR_U48 ( .A(R2_n1402), .Z(R2_n1338) );
  BUF_X1 R2_SR_U47 ( .A(R2_n1403), .Z(R2_n1339) );
  BUF_X1 R2_SR_U46 ( .A(R2_n1404), .Z(R2_n1340) );
  BUF_X1 R2_SR_U45 ( .A(R2_n1405), .Z(R2_n1341) );
  BUF_X1 R2_SR_U44 ( .A(R2_n1406), .Z(R2_n1342) );
  BUF_X1 R2_SR_U43 ( .A(R2_n1407), .Z(R2_n1343) );
  BUF_X1 R2_SR_U42 ( .A(R2_n1408), .Z(R2_n1344) );
  BUF_X1 R2_SR_U41 ( .A(R2_n1409), .Z(R2_n1345) );
  BUF_X1 R2_SR_U40 ( .A(R2_n1442), .Z(R2_n1346) );
  BUF_X1 R2_SR_U39 ( .A(R2_n1443), .Z(R2_n1347) );
  BUF_X1 R2_SR_U38 ( .A(R2_n1444), .Z(R2_n1348) );
  BUF_X1 R2_SR_U37 ( .A(R2_n1445), .Z(R2_n1349) );
  BUF_X1 R2_SR_U36 ( .A(R2_n1446), .Z(R2_n1350) );
  BUF_X1 R2_SR_U35 ( .A(R2_n1447), .Z(R2_n1351) );
  BUF_X1 R2_SR_U34 ( .A(R2_n1448), .Z(R2_n1352) );
  BUF_X1 R2_SR_U33 ( .A(R2_n1449), .Z(R2_n1353) );
  BUF_X1 R2_SR_U32 ( .A(R2_n1482), .Z(R2_n1354) );
  BUF_X1 R2_SR_U31 ( .A(R2_n1483), .Z(R2_n1355) );
  BUF_X1 R2_SR_U30 ( .A(R2_n1484), .Z(R2_n1356) );
  BUF_X1 R2_SR_U29 ( .A(R2_n1485), .Z(R2_n1357) );
  BUF_X1 R2_SR_U28 ( .A(R2_n1486), .Z(R2_n1358) );
  BUF_X1 R2_SR_U27 ( .A(R2_n1487), .Z(R2_n1359) );
  BUF_X1 R2_SR_U26 ( .A(R2_n1488), .Z(R2_n1360) );
  BUF_X1 R2_SR_U25 ( .A(R2_n1489), .Z(R2_n1361) );
  BUF_X1 R2_SR_U24 ( .A(R2_n1394), .Z(R2_n1362) );
  BUF_X1 R2_SR_U23 ( .A(R2_n1395), .Z(R2_n1363) );
  BUF_X1 R2_SR_U22 ( .A(R2_n1396), .Z(R2_n1364) );
  BUF_X1 R2_SR_U21 ( .A(R2_n1397), .Z(R2_n1365) );
  BUF_X1 R2_SR_U20 ( .A(R2_n1398), .Z(R2_n1366) );
  BUF_X1 R2_SR_U19 ( .A(R2_n1399), .Z(R2_n1367) );
  BUF_X1 R2_SR_U18 ( .A(R2_n1400), .Z(R2_n1368) );
  BUF_X1 R2_SR_U17 ( .A(R2_n1401), .Z(R2_n1369) );
  BUF_X1 R2_SR_U16 ( .A(R2_n1434), .Z(R2_n1370) );
  BUF_X1 R2_SR_U15 ( .A(R2_n1435), .Z(R2_n1371) );
  BUF_X1 R2_SR_U14 ( .A(R2_n1436), .Z(R2_n1372) );
  BUF_X1 R2_SR_U13 ( .A(R2_n1437), .Z(R2_n1373) );
  BUF_X1 R2_SR_U12 ( .A(R2_n1438), .Z(R2_n1374) );
  BUF_X1 R2_SR_U11 ( .A(R2_n1439), .Z(R2_n1375) );
  BUF_X1 R2_SR_U10 ( .A(R2_n1440), .Z(R2_n1376) );
  BUF_X1 R2_SR_U9 ( .A(R2_n1441), .Z(R2_n1377) );
  BUF_X1 R2_SR_U8 ( .A(R2_n1474), .Z(R2_n1378) );
  BUF_X1 R2_SR_U7 ( .A(R2_n1475), .Z(R2_n1379) );
  BUF_X1 R2_SR_U6 ( .A(R2_n1476), .Z(R2_n1380) );
  BUF_X1 R2_SR_U5 ( .A(R2_n1477), .Z(R2_n1381) );
  BUF_X1 R2_SR_U4 ( .A(R2_n1478), .Z(R2_n1382) );
  BUF_X1 R2_SR_U3 ( .A(R2_n1479), .Z(R2_n1383) );
  BUF_X1 R2_SR_U2 ( .A(R2_n1480), .Z(R2_n1384) );
  BUF_X1 R2_SR_U1 ( .A(R2_n1481), .Z(R2_n1385) );
  INV_X1 R2_MC1_U33 ( .A(R2_n1232), .ZN(R2_MC1_n4) );
  XOR2_X1 R2_MC1_U32 ( .A(R2_n1180), .B(R2_n1184), .Z(R2_MC1_n166) );
  XOR2_X1 R2_MC1_U31 ( .A(R2_n1212), .B(R2_n1216), .Z(R2_MC1_n76) );
  XNOR2_X1 R2_MC1_U30 ( .A(R2_n1225), .B(R2_MC1_n4), .ZN(R2_MC1_n31) );
  XNOR2_X1 R2_MC1_U29 ( .A(R2_n1228), .B(R2_MC1_n4), .ZN(R2_MC1_n280) );
  XNOR2_X1 R2_MC1_U28 ( .A(R2_n1172), .B(R2_MC1_n213), .ZN(R2_MC1_n146) );
  XNOR2_X1 R2_MC1_U27 ( .A(R2_n1204), .B(R2_MC1_n120), .ZN(R2_MC1_n53) );
  XNOR2_X1 R2_MC1_U26 ( .A(R2_n1180), .B(R2_n1164), .ZN(R2_MC1_n145) );
  XNOR2_X1 R2_MC1_U25 ( .A(R2_n1212), .B(R2_n1196), .ZN(R2_MC1_n52) );
  XOR2_X1 R2_MC1_U24 ( .A(R2_n1148), .B(R2_n1132), .Z(R2_MC1_n233) );
  XOR2_X1 R2_MC1_U23 ( .A(R2_n1244), .B(R2_n1228), .Z(R2_MC1_n283) );
  XNOR2_X1 R2_MC1_U22 ( .A(R2_n1236), .B(R2_MC1_n284), .ZN(R2_MC1_n23) );
  XNOR2_X1 R2_MC1_U21 ( .A(R2_n1140), .B(R2_MC1_n234), .ZN(R2_MC1_n201) );
  XNOR2_X1 R2_MC1_U20 ( .A(R2_n1171), .B(R2_n1176), .ZN(R2_MC1_n188) );
  XNOR2_X1 R2_MC1_U19 ( .A(R2_n1203), .B(R2_n1208), .ZN(R2_MC1_n96) );
  XNOR2_X1 R2_MC1_U18 ( .A(R2_n1155), .B(R2_n1160), .ZN(R2_MC1_n235) );
  XNOR2_X1 R2_MC1_U17 ( .A(R2_n1251), .B(R2_n1256), .ZN(R2_MC1_n285) );
  XNOR2_X1 R2_MC1_U16 ( .A(R2_n1172), .B(R2_n1164), .ZN(R2_MC1_n167) );
  INV_X1 R2_MC1_U15 ( .A(R2_MC1_n146), .ZN(R2_MC1_n11) );
  XNOR2_X1 R2_MC1_U14 ( .A(R2_MC1_n23), .B(R2_MC1_n24), .ZN(R2_MC1_n22) );
  XNOR2_X1 R2_MC1_U13 ( .A(R2_n1236), .B(R2_n1228), .ZN(R2_MC1_n306) );
  INV_X1 R2_MC1_U12 ( .A(R2_MC1_n285), .ZN(R2_MC1_n1) );
  XNOR2_X1 R2_MC1_U11 ( .A(R2_MC1_n201), .B(R2_MC1_n202), .ZN(R2_MC1_n200) );
  XNOR2_X1 R2_MC1_U10 ( .A(R2_n1140), .B(R2_n1132), .ZN(R2_MC1_n256) );
  INV_X1 R2_MC1_U9 ( .A(R2_MC1_n235), .ZN(R2_MC1_n13) );
  XNOR2_X1 R2_MC1_U8 ( .A(R2_n1204), .B(R2_n1196), .ZN(R2_MC1_n77) );
  INV_X1 R2_MC1_U7 ( .A(R2_MC1_n53), .ZN(R2_MC1_n7) );
  XNOR2_X1 R2_MC1_U6 ( .A(R2_MC1_n201), .B(R2_MC1_n233), .ZN(R2_MC1_n232) );
  XNOR2_X1 R2_MC1_U5 ( .A(R2_MC1_n144), .B(R2_MC1_n169), .ZN(R2_MC1_n168) );
  XNOR2_X1 R2_MC1_U4 ( .A(R2_MC1_n51), .B(R2_MC1_n79), .ZN(R2_MC1_n78) );
  XNOR2_X1 R2_MC1_U3 ( .A(R2_MC1_n23), .B(R2_MC1_n283), .ZN(R2_MC1_n282) );
  XNOR2_X1 R2_MC1_U2 ( .A(R2_MC1_n145), .B(R2_MC1_n144), .ZN(R2_MC1_n143) );
  XNOR2_X1 R2_MC1_U1 ( .A(R2_MC1_n52), .B(R2_MC1_n51), .ZN(R2_MC1_n50) );
  XOR2_X1 R2_MC1_U466 ( .A(R2_n1144), .B(R2_n1136), .Z(R2_MC1_n219) );
  XOR2_X1 R2_MC1_U465 ( .A(R2_n1153), .B(R2_n1145), .Z(R2_MC1_n59) );
  XOR2_X1 R2_MC1_U464 ( .A(R2_n1137), .B(R2_MC1_n59), .Z(R2_MC1_n338) );
  XOR2_X1 R2_MC1_U463 ( .A(R2_MC1_n219), .B(R2_MC1_n338), .Z(R2_U16_DATA2_0)
         );
  XOR2_X1 R2_MC1_U462 ( .A(R2_n1237), .B(R2_n1245), .Z(R2_MC1_n279) );
  XOR2_X1 R2_MC1_U461 ( .A(R2_n1253), .B(R2_MC1_n279), .Z(R2_MC1_n336) );
  XOR2_X1 R2_MC1_U460 ( .A(R2_n1236), .B(R2_n1240), .Z(R2_MC1_n322) );
  XOR2_X1 R2_MC1_U459 ( .A(R2_MC1_n280), .B(R2_MC1_n322), .Z(R2_MC1_n337) );
  XOR2_X1 R2_MC1_U458 ( .A(R2_MC1_n336), .B(R2_MC1_n337), .Z(R2_U16_DATA2_100)
         );
  XOR2_X1 R2_MC1_U457 ( .A(R2_n1254), .B(R2_n1237), .Z(R2_MC1_n334) );
  XOR2_X1 R2_MC1_U456 ( .A(R2_n1238), .B(R2_n1246), .Z(R2_MC1_n274) );
  XOR2_X1 R2_MC1_U455 ( .A(R2_n1229), .B(R2_MC1_n274), .Z(R2_MC1_n335) );
  XOR2_X1 R2_MC1_U454 ( .A(R2_MC1_n334), .B(R2_MC1_n335), .Z(R2_U16_DATA2_101)
         );
  XOR2_X1 R2_MC1_U453 ( .A(R2_n1255), .B(R2_n1238), .Z(R2_MC1_n332) );
  XOR2_X1 R2_MC1_U452 ( .A(R2_n1239), .B(R2_n1247), .Z(R2_MC1_n271) );
  XOR2_X1 R2_MC1_U451 ( .A(R2_n1230), .B(R2_MC1_n271), .Z(R2_MC1_n333) );
  XOR2_X1 R2_MC1_U450 ( .A(R2_MC1_n332), .B(R2_MC1_n333), .Z(R2_U16_DATA2_102)
         );
  XOR2_X1 R2_MC1_U449 ( .A(R2_n1240), .B(R2_n1239), .Z(R2_MC1_n330) );
  XOR2_X1 R2_MC1_U448 ( .A(R2_n1248), .B(R2_n1256), .Z(R2_MC1_n314) );
  XOR2_X1 R2_MC1_U447 ( .A(R2_n1231), .B(R2_MC1_n314), .Z(R2_MC1_n331) );
  XOR2_X1 R2_MC1_U446 ( .A(R2_MC1_n330), .B(R2_MC1_n331), .Z(R2_U16_DATA2_103)
         );
  XOR2_X1 R2_MC1_U445 ( .A(R2_n1248), .B(R2_n1240), .Z(R2_MC1_n328) );
  XOR2_X1 R2_MC1_U444 ( .A(R2_n1249), .B(R2_n1241), .Z(R2_MC1_n35) );
  XOR2_X1 R2_MC1_U443 ( .A(R2_n1225), .B(R2_MC1_n35), .Z(R2_MC1_n329) );
  XOR2_X1 R2_MC1_U442 ( .A(R2_MC1_n328), .B(R2_MC1_n329), .Z(R2_U16_DATA2_104)
         );
  XOR2_X1 R2_MC1_U441 ( .A(R2_n1233), .B(R2_n1240), .Z(R2_MC1_n30) );
  XOR2_X1 R2_MC1_U440 ( .A(R2_n1242), .B(R2_MC1_n30), .Z(R2_MC1_n326) );
  XOR2_X1 R2_MC1_U439 ( .A(R2_n1250), .B(R2_n1226), .Z(R2_MC1_n286) );
  XOR2_X1 R2_MC1_U438 ( .A(R2_n1241), .B(R2_n1248), .Z(R2_MC1_n313) );
  XOR2_X1 R2_MC1_U437 ( .A(R2_MC1_n286), .B(R2_MC1_n313), .Z(R2_MC1_n327) );
  XOR2_X1 R2_MC1_U436 ( .A(R2_MC1_n326), .B(R2_MC1_n327), .Z(R2_U16_DATA2_105)
         );
  XOR2_X1 R2_MC1_U435 ( .A(R2_n1234), .B(R2_n1242), .Z(R2_MC1_n32) );
  XOR2_X1 R2_MC1_U434 ( .A(R2_n1251), .B(R2_n1243), .Z(R2_MC1_n27) );
  XOR2_X1 R2_MC1_U433 ( .A(R2_n1227), .B(R2_MC1_n27), .Z(R2_MC1_n325) );
  XOR2_X1 R2_MC1_U432 ( .A(R2_MC1_n32), .B(R2_MC1_n325), .Z(R2_U16_DATA2_106)
         );
  XOR2_X1 R2_MC1_U431 ( .A(R2_n1248), .B(R2_n1243), .Z(R2_MC1_n324) );
  XOR2_X1 R2_MC1_U430 ( .A(R2_n1252), .B(R2_MC1_n324), .Z(R2_MC1_n308) );
  XOR2_X1 R2_MC1_U429 ( .A(R2_n1235), .B(R2_n1240), .Z(R2_MC1_n24) );
  XOR2_X1 R2_MC1_U428 ( .A(R2_MC1_n24), .B(R2_MC1_n283), .Z(R2_MC1_n323) );
  XOR2_X1 R2_MC1_U427 ( .A(R2_MC1_n308), .B(R2_MC1_n323), .Z(R2_U16_DATA2_107)
         );
  XOR2_X1 R2_MC1_U426 ( .A(R2_n1229), .B(R2_n1253), .Z(R2_MC1_n276) );
  XOR2_X1 R2_MC1_U425 ( .A(R2_n1245), .B(R2_MC1_n276), .Z(R2_MC1_n320) );
  XOR2_X1 R2_MC1_U424 ( .A(R2_n1244), .B(R2_n1248), .Z(R2_MC1_n305) );
  XOR2_X1 R2_MC1_U423 ( .A(R2_MC1_n305), .B(R2_MC1_n322), .Z(R2_MC1_n321) );
  XOR2_X1 R2_MC1_U422 ( .A(R2_MC1_n320), .B(R2_MC1_n321), .Z(R2_U16_DATA2_108)
         );
  XOR2_X1 R2_MC1_U421 ( .A(R2_n1230), .B(R2_n1254), .Z(R2_MC1_n273) );
  XOR2_X1 R2_MC1_U420 ( .A(R2_n1246), .B(R2_MC1_n273), .Z(R2_MC1_n319) );
  XOR2_X1 R2_MC1_U419 ( .A(R2_MC1_n279), .B(R2_MC1_n319), .Z(R2_U16_DATA2_109)
         );
  XOR2_X1 R2_MC1_U418 ( .A(R2_n1146), .B(R2_n1138), .Z(R2_MC1_n254) );
  XOR2_X1 R2_MC1_U417 ( .A(R2_n1155), .B(R2_n1147), .Z(R2_MC1_n226) );
  XOR2_X1 R2_MC1_U416 ( .A(R2_n1131), .B(R2_MC1_n226), .Z(R2_MC1_n318) );
  XOR2_X1 R2_MC1_U415 ( .A(R2_MC1_n254), .B(R2_MC1_n318), .Z(R2_U16_DATA2_10)
         );
  XOR2_X1 R2_MC1_U414 ( .A(R2_n1231), .B(R2_n1255), .Z(R2_MC1_n269) );
  XOR2_X1 R2_MC1_U413 ( .A(R2_n1247), .B(R2_MC1_n269), .Z(R2_MC1_n317) );
  XOR2_X1 R2_MC1_U412 ( .A(R2_MC1_n274), .B(R2_MC1_n317), .Z(R2_U16_DATA2_110)
         );
  XOR2_X1 R2_MC1_U411 ( .A(R2_n1232), .B(R2_MC1_n271), .Z(R2_MC1_n316) );
  XOR2_X1 R2_MC1_U410 ( .A(R2_MC1_n314), .B(R2_MC1_n316), .Z(R2_U16_DATA2_111)
         );
  XOR2_X1 R2_MC1_U409 ( .A(R2_n1233), .B(R2_n1225), .Z(R2_MC1_n294) );
  XOR2_X1 R2_MC1_U408 ( .A(R2_n1249), .B(R2_MC1_n294), .Z(R2_MC1_n315) );
  XOR2_X1 R2_MC1_U407 ( .A(R2_MC1_n314), .B(R2_MC1_n315), .Z(R2_U16_DATA2_112)
         );
  XOR2_X1 R2_MC1_U406 ( .A(R2_n1234), .B(R2_MC1_n286), .Z(R2_MC1_n311) );
  XOR2_X1 R2_MC1_U405 ( .A(R2_n1249), .B(R2_n1256), .Z(R2_MC1_n291) );
  XOR2_X1 R2_MC1_U404 ( .A(R2_MC1_n291), .B(R2_MC1_n313), .Z(R2_MC1_n312) );
  XOR2_X1 R2_MC1_U403 ( .A(R2_MC1_n311), .B(R2_MC1_n312), .Z(R2_U16_DATA2_113)
         );
  XOR2_X1 R2_MC1_U402 ( .A(R2_n1250), .B(R2_n1242), .Z(R2_MC1_n309) );
  XOR2_X1 R2_MC1_U401 ( .A(R2_n1235), .B(R2_n1227), .Z(R2_MC1_n288) );
  XOR2_X1 R2_MC1_U400 ( .A(R2_n1251), .B(R2_MC1_n288), .Z(R2_MC1_n310) );
  XOR2_X1 R2_MC1_U399 ( .A(R2_MC1_n309), .B(R2_MC1_n310), .Z(R2_U16_DATA2_114)
         );
  XOR2_X1 R2_MC1_U397 ( .A(R2_MC1_n285), .B(R2_MC1_n308), .Z(R2_MC1_n307) );
  XOR2_X1 R2_MC1_U396 ( .A(R2_MC1_n306), .B(R2_MC1_n307), .Z(R2_U16_DATA2_115)
         );
  XOR2_X1 R2_MC1_U395 ( .A(R2_n1237), .B(R2_MC1_n276), .Z(R2_MC1_n303) );
  XOR2_X1 R2_MC1_U394 ( .A(R2_n1252), .B(R2_n1256), .Z(R2_MC1_n281) );
  XOR2_X1 R2_MC1_U393 ( .A(R2_MC1_n281), .B(R2_MC1_n305), .Z(R2_MC1_n304) );
  XOR2_X1 R2_MC1_U392 ( .A(R2_MC1_n303), .B(R2_MC1_n304), .Z(R2_U16_DATA2_116)
         );
  XOR2_X1 R2_MC1_U391 ( .A(R2_n1253), .B(R2_n1245), .Z(R2_MC1_n301) );
  XOR2_X1 R2_MC1_U390 ( .A(R2_n1238), .B(R2_MC1_n273), .Z(R2_MC1_n302) );
  XOR2_X1 R2_MC1_U389 ( .A(R2_MC1_n301), .B(R2_MC1_n302), .Z(R2_U16_DATA2_117)
         );
  XOR2_X1 R2_MC1_U388 ( .A(R2_n1254), .B(R2_n1246), .Z(R2_MC1_n299) );
  XOR2_X1 R2_MC1_U387 ( .A(R2_n1239), .B(R2_MC1_n269), .Z(R2_MC1_n300) );
  XOR2_X1 R2_MC1_U386 ( .A(R2_MC1_n299), .B(R2_MC1_n300), .Z(R2_U16_DATA2_118)
         );
  XOR2_X1 R2_MC1_U385 ( .A(R2_n1256), .B(R2_n1255), .Z(R2_MC1_n297) );
  XOR2_X1 R2_MC1_U384 ( .A(R2_n1232), .B(R2_n1240), .Z(R2_MC1_n33) );
  XOR2_X1 R2_MC1_U383 ( .A(R2_n1247), .B(R2_MC1_n33), .Z(R2_MC1_n298) );
  XOR2_X1 R2_MC1_U382 ( .A(R2_MC1_n297), .B(R2_MC1_n298), .Z(R2_U16_DATA2_119)
         );
  XOR2_X1 R2_MC1_U381 ( .A(R2_n1152), .B(R2_n1147), .Z(R2_MC1_n296) );
  XOR2_X1 R2_MC1_U380 ( .A(R2_n1156), .B(R2_MC1_n296), .Z(R2_MC1_n258) );
  XOR2_X1 R2_MC1_U379 ( .A(R2_n1139), .B(R2_n1144), .Z(R2_MC1_n202) );
  XOR2_X1 R2_MC1_U378 ( .A(R2_MC1_n202), .B(R2_MC1_n233), .Z(R2_MC1_n295) );
  XOR2_X1 R2_MC1_U377 ( .A(R2_MC1_n258), .B(R2_MC1_n295), .Z(R2_U16_DATA2_11)
         );
  XOR2_X1 R2_MC1_U376 ( .A(R2_n1256), .B(R2_n1232), .Z(R2_MC1_n292) );
  XOR2_X1 R2_MC1_U375 ( .A(R2_n1241), .B(R2_MC1_n294), .Z(R2_MC1_n293) );
  XOR2_X1 R2_MC1_U374 ( .A(R2_MC1_n292), .B(R2_MC1_n293), .Z(R2_U16_DATA2_120)
         );
  XOR2_X1 R2_MC1_U373 ( .A(R2_n1226), .B(R2_MC1_n32), .Z(R2_MC1_n289) );
  XOR2_X1 R2_MC1_U372 ( .A(R2_MC1_n31), .B(R2_MC1_n291), .Z(R2_MC1_n290) );
  XOR2_X1 R2_MC1_U371 ( .A(R2_MC1_n289), .B(R2_MC1_n290), .Z(R2_U16_DATA2_121)
         );
  XOR2_X1 R2_MC1_U370 ( .A(R2_n1243), .B(R2_MC1_n288), .Z(R2_MC1_n287) );
  XOR2_X1 R2_MC1_U369 ( .A(R2_MC1_n286), .B(R2_MC1_n287), .Z(R2_U16_DATA2_122)
         );
  XOR2_X1 R2_MC1_U368 ( .A(R2_n1232), .B(R2_n1227), .Z(R2_MC1_n284) );
  XOR2_X1 R2_MC1_U367 ( .A(R2_MC1_n1), .B(R2_MC1_n282), .Z(R2_U16_DATA2_123)
         );
  XOR2_X1 R2_MC1_U366 ( .A(R2_n1229), .B(R2_MC1_n281), .Z(R2_MC1_n277) );
  XOR2_X1 R2_MC1_U365 ( .A(R2_MC1_n279), .B(R2_MC1_n280), .Z(R2_MC1_n278) );
  XOR2_X1 R2_MC1_U364 ( .A(R2_MC1_n277), .B(R2_MC1_n278), .Z(R2_U16_DATA2_124)
         );
  XOR2_X1 R2_MC1_U363 ( .A(R2_n1230), .B(R2_MC1_n276), .Z(R2_MC1_n275) );
  XOR2_X1 R2_MC1_U362 ( .A(R2_MC1_n274), .B(R2_MC1_n275), .Z(R2_U16_DATA2_125)
         );
  XOR2_X1 R2_MC1_U361 ( .A(R2_n1231), .B(R2_MC1_n273), .Z(R2_MC1_n272) );
  XOR2_X1 R2_MC1_U360 ( .A(R2_MC1_n271), .B(R2_MC1_n272), .Z(R2_U16_DATA2_126)
         );
  XOR2_X1 R2_MC1_U359 ( .A(R2_n1248), .B(R2_MC1_n33), .Z(R2_MC1_n270) );
  XOR2_X1 R2_MC1_U358 ( .A(R2_MC1_n269), .B(R2_MC1_n270), .Z(R2_U16_DATA2_127)
         );
  XOR2_X1 R2_MC1_U357 ( .A(R2_n1140), .B(R2_n1144), .Z(R2_MC1_n175) );
  XOR2_X1 R2_MC1_U356 ( .A(R2_n1149), .B(R2_MC1_n175), .Z(R2_MC1_n267) );
  XOR2_X1 R2_MC1_U355 ( .A(R2_n1157), .B(R2_n1133), .Z(R2_MC1_n227) );
  XOR2_X1 R2_MC1_U354 ( .A(R2_n1148), .B(R2_n1152), .Z(R2_MC1_n252) );
  XOR2_X1 R2_MC1_U353 ( .A(R2_MC1_n227), .B(R2_MC1_n252), .Z(R2_MC1_n268) );
  XOR2_X1 R2_MC1_U352 ( .A(R2_MC1_n267), .B(R2_MC1_n268), .Z(R2_U16_DATA2_12)
         );
  XOR2_X1 R2_MC1_U351 ( .A(R2_n1158), .B(R2_n1134), .Z(R2_MC1_n222) );
  XOR2_X1 R2_MC1_U350 ( .A(R2_n1141), .B(R2_n1149), .Z(R2_MC1_n176) );
  XOR2_X1 R2_MC1_U349 ( .A(R2_n1150), .B(R2_MC1_n176), .Z(R2_MC1_n266) );
  XOR2_X1 R2_MC1_U348 ( .A(R2_MC1_n222), .B(R2_MC1_n266), .Z(R2_U16_DATA2_13)
         );
  XOR2_X1 R2_MC1_U347 ( .A(R2_n1159), .B(R2_n1135), .Z(R2_MC1_n221) );
  XOR2_X1 R2_MC1_U346 ( .A(R2_n1142), .B(R2_n1150), .Z(R2_MC1_n142) );
  XOR2_X1 R2_MC1_U345 ( .A(R2_n1151), .B(R2_MC1_n142), .Z(R2_MC1_n265) );
  XOR2_X1 R2_MC1_U344 ( .A(R2_MC1_n221), .B(R2_MC1_n265), .Z(R2_U16_DATA2_14)
         );
  XOR2_X1 R2_MC1_U343 ( .A(R2_n1143), .B(R2_n1151), .Z(R2_MC1_n113) );
  XOR2_X1 R2_MC1_U342 ( .A(R2_n1152), .B(R2_n1160), .Z(R2_MC1_n89) );
  XOR2_X1 R2_MC1_U341 ( .A(R2_n1136), .B(R2_MC1_n89), .Z(R2_MC1_n264) );
  XOR2_X1 R2_MC1_U340 ( .A(R2_MC1_n113), .B(R2_MC1_n264), .Z(R2_U16_DATA2_15)
         );
  XOR2_X1 R2_MC1_U339 ( .A(R2_n1137), .B(R2_n1129), .Z(R2_MC1_n243) );
  XOR2_X1 R2_MC1_U338 ( .A(R2_n1153), .B(R2_MC1_n89), .Z(R2_MC1_n263) );
  XOR2_X1 R2_MC1_U337 ( .A(R2_MC1_n243), .B(R2_MC1_n263), .Z(R2_U16_DATA2_16)
         );
  XOR2_X1 R2_MC1_U336 ( .A(R2_n1130), .B(R2_n1154), .Z(R2_MC1_n20) );
  XOR2_X1 R2_MC1_U335 ( .A(R2_n1138), .B(R2_MC1_n20), .Z(R2_MC1_n261) );
  XOR2_X1 R2_MC1_U334 ( .A(R2_n1145), .B(R2_n1152), .Z(R2_MC1_n18) );
  XOR2_X1 R2_MC1_U333 ( .A(R2_n1153), .B(R2_n1160), .Z(R2_MC1_n240) );
  XOR2_X1 R2_MC1_U332 ( .A(R2_MC1_n18), .B(R2_MC1_n240), .Z(R2_MC1_n262) );
  XOR2_X1 R2_MC1_U331 ( .A(R2_MC1_n261), .B(R2_MC1_n262), .Z(R2_U16_DATA2_17)
         );
  XOR2_X1 R2_MC1_U330 ( .A(R2_n1154), .B(R2_n1146), .Z(R2_MC1_n259) );
  XOR2_X1 R2_MC1_U329 ( .A(R2_n1139), .B(R2_n1131), .Z(R2_MC1_n236) );
  XOR2_X1 R2_MC1_U328 ( .A(R2_n1155), .B(R2_MC1_n236), .Z(R2_MC1_n260) );
  XOR2_X1 R2_MC1_U327 ( .A(R2_MC1_n259), .B(R2_MC1_n260), .Z(R2_U16_DATA2_18)
         );
  XOR2_X1 R2_MC1_U325 ( .A(R2_MC1_n235), .B(R2_MC1_n258), .Z(R2_MC1_n257) );
  XOR2_X1 R2_MC1_U324 ( .A(R2_MC1_n256), .B(R2_MC1_n257), .Z(R2_U16_DATA2_19)
         );
  XOR2_X1 R2_MC1_U323 ( .A(R2_n1137), .B(R2_n1144), .Z(R2_MC1_n19) );
  XOR2_X1 R2_MC1_U322 ( .A(R2_n1154), .B(R2_MC1_n19), .Z(R2_MC1_n253) );
  XOR2_X1 R2_MC1_U321 ( .A(R2_n1129), .B(R2_n1136), .Z(R2_MC1_n255) );
  XOR2_X1 R2_MC1_U320 ( .A(R2_MC1_n254), .B(R2_MC1_n255), .Z(R2_MC1_n239) );
  XOR2_X1 R2_MC1_U319 ( .A(R2_MC1_n253), .B(R2_MC1_n239), .Z(R2_U16_DATA2_1)
         );
  XOR2_X1 R2_MC1_U318 ( .A(R2_n1141), .B(R2_MC1_n227), .Z(R2_MC1_n250) );
  XOR2_X1 R2_MC1_U317 ( .A(R2_n1156), .B(R2_n1160), .Z(R2_MC1_n231) );
  XOR2_X1 R2_MC1_U316 ( .A(R2_MC1_n231), .B(R2_MC1_n252), .Z(R2_MC1_n251) );
  XOR2_X1 R2_MC1_U315 ( .A(R2_MC1_n250), .B(R2_MC1_n251), .Z(R2_U16_DATA2_20)
         );
  XOR2_X1 R2_MC1_U314 ( .A(R2_n1157), .B(R2_n1149), .Z(R2_MC1_n248) );
  XOR2_X1 R2_MC1_U313 ( .A(R2_n1142), .B(R2_MC1_n222), .Z(R2_MC1_n249) );
  XOR2_X1 R2_MC1_U312 ( .A(R2_MC1_n248), .B(R2_MC1_n249), .Z(R2_U16_DATA2_21)
         );
  XOR2_X1 R2_MC1_U311 ( .A(R2_n1158), .B(R2_n1150), .Z(R2_MC1_n246) );
  XOR2_X1 R2_MC1_U310 ( .A(R2_n1143), .B(R2_MC1_n221), .Z(R2_MC1_n247) );
  XOR2_X1 R2_MC1_U309 ( .A(R2_MC1_n246), .B(R2_MC1_n247), .Z(R2_U16_DATA2_22)
         );
  XOR2_X1 R2_MC1_U308 ( .A(R2_n1160), .B(R2_n1159), .Z(R2_MC1_n244) );
  XOR2_X1 R2_MC1_U307 ( .A(R2_n1151), .B(R2_MC1_n219), .Z(R2_MC1_n245) );
  XOR2_X1 R2_MC1_U306 ( .A(R2_MC1_n244), .B(R2_MC1_n245), .Z(R2_U16_DATA2_23)
         );
  XOR2_X1 R2_MC1_U305 ( .A(R2_n1136), .B(R2_n1160), .Z(R2_MC1_n241) );
  XOR2_X1 R2_MC1_U304 ( .A(R2_n1145), .B(R2_MC1_n243), .Z(R2_MC1_n242) );
  XOR2_X1 R2_MC1_U303 ( .A(R2_MC1_n241), .B(R2_MC1_n242), .Z(R2_U16_DATA2_24)
         );
  XOR2_X1 R2_MC1_U302 ( .A(R2_n1130), .B(R2_MC1_n240), .Z(R2_MC1_n238) );
  XOR2_X1 R2_MC1_U301 ( .A(R2_MC1_n238), .B(R2_MC1_n239), .Z(R2_U16_DATA2_25)
         );
  XOR2_X1 R2_MC1_U300 ( .A(R2_n1147), .B(R2_MC1_n20), .Z(R2_MC1_n237) );
  XOR2_X1 R2_MC1_U299 ( .A(R2_MC1_n236), .B(R2_MC1_n237), .Z(R2_U16_DATA2_26)
         );
  XOR2_X1 R2_MC1_U298 ( .A(R2_n1136), .B(R2_n1131), .Z(R2_MC1_n234) );
  XOR2_X1 R2_MC1_U297 ( .A(R2_MC1_n13), .B(R2_MC1_n232), .Z(R2_U16_DATA2_27)
         );
  XOR2_X1 R2_MC1_U296 ( .A(R2_n1133), .B(R2_MC1_n176), .Z(R2_MC1_n229) );
  XOR2_X1 R2_MC1_U295 ( .A(R2_n1132), .B(R2_n1136), .Z(R2_MC1_n174) );
  XOR2_X1 R2_MC1_U294 ( .A(R2_MC1_n174), .B(R2_MC1_n231), .Z(R2_MC1_n230) );
  XOR2_X1 R2_MC1_U293 ( .A(R2_MC1_n229), .B(R2_MC1_n230), .Z(R2_U16_DATA2_28)
         );
  XOR2_X1 R2_MC1_U292 ( .A(R2_n1134), .B(R2_MC1_n142), .Z(R2_MC1_n228) );
  XOR2_X1 R2_MC1_U291 ( .A(R2_MC1_n227), .B(R2_MC1_n228), .Z(R2_U16_DATA2_29)
         );
  XOR2_X1 R2_MC1_U290 ( .A(R2_n1138), .B(R2_n1130), .Z(R2_MC1_n224) );
  XOR2_X1 R2_MC1_U289 ( .A(R2_n1139), .B(R2_MC1_n226), .Z(R2_MC1_n225) );
  XOR2_X1 R2_MC1_U288 ( .A(R2_MC1_n224), .B(R2_MC1_n225), .Z(R2_U16_DATA2_2)
         );
  XOR2_X1 R2_MC1_U287 ( .A(R2_n1135), .B(R2_MC1_n113), .Z(R2_MC1_n223) );
  XOR2_X1 R2_MC1_U286 ( .A(R2_MC1_n222), .B(R2_MC1_n223), .Z(R2_U16_DATA2_30)
         );
  XOR2_X1 R2_MC1_U285 ( .A(R2_n1152), .B(R2_MC1_n221), .Z(R2_MC1_n220) );
  XOR2_X1 R2_MC1_U284 ( .A(R2_MC1_n219), .B(R2_MC1_n220), .Z(R2_U16_DATA2_31)
         );
  XOR2_X1 R2_MC1_U283 ( .A(R2_n1185), .B(R2_n1177), .Z(R2_MC1_n198) );
  XOR2_X1 R2_MC1_U282 ( .A(R2_n1168), .B(R2_n1176), .Z(R2_MC1_n126) );
  XOR2_X1 R2_MC1_U281 ( .A(R2_n1169), .B(R2_MC1_n126), .Z(R2_MC1_n218) );
  XOR2_X1 R2_MC1_U280 ( .A(R2_MC1_n198), .B(R2_MC1_n218), .Z(R2_U16_DATA2_32)
         );
  XOR2_X1 R2_MC1_U279 ( .A(R2_n1170), .B(R2_n1178), .Z(R2_MC1_n152) );
  XOR2_X1 R2_MC1_U278 ( .A(R2_n1186), .B(R2_MC1_n152), .Z(R2_MC1_n216) );
  XOR2_X1 R2_MC1_U277 ( .A(R2_n1161), .B(R2_n1168), .Z(R2_MC1_n153) );
  XOR2_X1 R2_MC1_U276 ( .A(R2_n1169), .B(R2_n1176), .Z(R2_MC1_n195) );
  XOR2_X1 R2_MC1_U275 ( .A(R2_MC1_n153), .B(R2_MC1_n195), .Z(R2_MC1_n217) );
  XOR2_X1 R2_MC1_U274 ( .A(R2_MC1_n216), .B(R2_MC1_n217), .Z(R2_U16_DATA2_33)
         );
  XOR2_X1 R2_MC1_U273 ( .A(R2_n1170), .B(R2_n1162), .Z(R2_MC1_n214) );
  XOR2_X1 R2_MC1_U272 ( .A(R2_n1187), .B(R2_n1179), .Z(R2_MC1_n191) );
  XOR2_X1 R2_MC1_U271 ( .A(R2_n1171), .B(R2_MC1_n191), .Z(R2_MC1_n215) );
  XOR2_X1 R2_MC1_U270 ( .A(R2_MC1_n214), .B(R2_MC1_n215), .Z(R2_U16_DATA2_34)
         );
  XOR2_X1 R2_MC1_U269 ( .A(R2_n1180), .B(R2_n1188), .Z(R2_MC1_n211) );
  XOR2_X1 R2_MC1_U268 ( .A(R2_n1168), .B(R2_n1163), .Z(R2_MC1_n213) );
  XOR2_X1 R2_MC1_U266 ( .A(R2_MC1_n146), .B(R2_MC1_n188), .Z(R2_MC1_n212) );
  XOR2_X1 R2_MC1_U265 ( .A(R2_MC1_n211), .B(R2_MC1_n212), .Z(R2_U16_DATA2_35)
         );
  XOR2_X1 R2_MC1_U264 ( .A(R2_n1173), .B(R2_n1181), .Z(R2_MC1_n137) );
  XOR2_X1 R2_MC1_U263 ( .A(R2_n1189), .B(R2_MC1_n137), .Z(R2_MC1_n209) );
  XOR2_X1 R2_MC1_U262 ( .A(R2_n1164), .B(R2_n1168), .Z(R2_MC1_n138) );
  XOR2_X1 R2_MC1_U261 ( .A(R2_n1172), .B(R2_n1176), .Z(R2_MC1_n187) );
  XOR2_X1 R2_MC1_U260 ( .A(R2_MC1_n138), .B(R2_MC1_n187), .Z(R2_MC1_n210) );
  XOR2_X1 R2_MC1_U259 ( .A(R2_MC1_n209), .B(R2_MC1_n210), .Z(R2_U16_DATA2_36)
         );
  XOR2_X1 R2_MC1_U258 ( .A(R2_n1190), .B(R2_n1173), .Z(R2_MC1_n207) );
  XOR2_X1 R2_MC1_U257 ( .A(R2_n1174), .B(R2_n1182), .Z(R2_MC1_n132) );
  XOR2_X1 R2_MC1_U256 ( .A(R2_n1165), .B(R2_MC1_n132), .Z(R2_MC1_n208) );
  XOR2_X1 R2_MC1_U255 ( .A(R2_MC1_n207), .B(R2_MC1_n208), .Z(R2_U16_DATA2_37)
         );
  XOR2_X1 R2_MC1_U254 ( .A(R2_n1191), .B(R2_n1174), .Z(R2_MC1_n205) );
  XOR2_X1 R2_MC1_U253 ( .A(R2_n1175), .B(R2_n1183), .Z(R2_MC1_n129) );
  XOR2_X1 R2_MC1_U252 ( .A(R2_n1166), .B(R2_MC1_n129), .Z(R2_MC1_n206) );
  XOR2_X1 R2_MC1_U251 ( .A(R2_MC1_n205), .B(R2_MC1_n206), .Z(R2_U16_DATA2_38)
         );
  XOR2_X1 R2_MC1_U250 ( .A(R2_n1176), .B(R2_n1175), .Z(R2_MC1_n203) );
  XOR2_X1 R2_MC1_U249 ( .A(R2_n1184), .B(R2_n1192), .Z(R2_MC1_n180) );
  XOR2_X1 R2_MC1_U248 ( .A(R2_n1167), .B(R2_MC1_n180), .Z(R2_MC1_n204) );
  XOR2_X1 R2_MC1_U247 ( .A(R2_MC1_n203), .B(R2_MC1_n204), .Z(R2_U16_DATA2_39)
         );
  XOR2_X1 R2_MC1_U246 ( .A(R2_n1148), .B(R2_n1156), .Z(R2_MC1_n199) );
  XOR2_X1 R2_MC1_U245 ( .A(R2_MC1_n199), .B(R2_MC1_n200), .Z(R2_U16_DATA2_3)
         );
  XOR2_X1 R2_MC1_U244 ( .A(R2_n1184), .B(R2_n1176), .Z(R2_MC1_n196) );
  XOR2_X1 R2_MC1_U243 ( .A(R2_n1161), .B(R2_MC1_n198), .Z(R2_MC1_n197) );
  XOR2_X1 R2_MC1_U242 ( .A(R2_MC1_n196), .B(R2_MC1_n197), .Z(R2_U16_DATA2_40)
         );
  XOR2_X1 R2_MC1_U241 ( .A(R2_n1162), .B(R2_n1186), .Z(R2_MC1_n147) );
  XOR2_X1 R2_MC1_U240 ( .A(R2_n1178), .B(R2_MC1_n147), .Z(R2_MC1_n193) );
  XOR2_X1 R2_MC1_U239 ( .A(R2_n1177), .B(R2_n1184), .Z(R2_MC1_n179) );
  XOR2_X1 R2_MC1_U238 ( .A(R2_MC1_n179), .B(R2_MC1_n195), .Z(R2_MC1_n194) );
  XOR2_X1 R2_MC1_U237 ( .A(R2_MC1_n193), .B(R2_MC1_n194), .Z(R2_U16_DATA2_41)
         );
  XOR2_X1 R2_MC1_U236 ( .A(R2_n1163), .B(R2_MC1_n152), .Z(R2_MC1_n192) );
  XOR2_X1 R2_MC1_U235 ( .A(R2_MC1_n191), .B(R2_MC1_n192), .Z(R2_U16_DATA2_42)
         );
  XOR2_X1 R2_MC1_U234 ( .A(R2_n1184), .B(R2_n1179), .Z(R2_MC1_n190) );
  XOR2_X1 R2_MC1_U233 ( .A(R2_n1188), .B(R2_MC1_n190), .Z(R2_MC1_n169) );
  XOR2_X1 R2_MC1_U232 ( .A(R2_MC1_n145), .B(R2_MC1_n169), .Z(R2_MC1_n189) );
  XOR2_X1 R2_MC1_U231 ( .A(R2_MC1_n188), .B(R2_MC1_n189), .Z(R2_U16_DATA2_43)
         );
  XOR2_X1 R2_MC1_U230 ( .A(R2_n1165), .B(R2_n1189), .Z(R2_MC1_n134) );
  XOR2_X1 R2_MC1_U229 ( .A(R2_n1181), .B(R2_MC1_n134), .Z(R2_MC1_n185) );
  XOR2_X1 R2_MC1_U228 ( .A(R2_MC1_n166), .B(R2_MC1_n187), .Z(R2_MC1_n186) );
  XOR2_X1 R2_MC1_U227 ( .A(R2_MC1_n185), .B(R2_MC1_n186), .Z(R2_U16_DATA2_44)
         );
  XOR2_X1 R2_MC1_U226 ( .A(R2_n1166), .B(R2_n1190), .Z(R2_MC1_n131) );
  XOR2_X1 R2_MC1_U225 ( .A(R2_n1182), .B(R2_MC1_n131), .Z(R2_MC1_n184) );
  XOR2_X1 R2_MC1_U224 ( .A(R2_MC1_n137), .B(R2_MC1_n184), .Z(R2_U16_DATA2_45)
         );
  XOR2_X1 R2_MC1_U223 ( .A(R2_n1167), .B(R2_n1191), .Z(R2_MC1_n128) );
  XOR2_X1 R2_MC1_U222 ( .A(R2_n1183), .B(R2_MC1_n128), .Z(R2_MC1_n183) );
  XOR2_X1 R2_MC1_U221 ( .A(R2_MC1_n132), .B(R2_MC1_n183), .Z(R2_U16_DATA2_46)
         );
  XOR2_X1 R2_MC1_U220 ( .A(R2_n1168), .B(R2_MC1_n129), .Z(R2_MC1_n182) );
  XOR2_X1 R2_MC1_U219 ( .A(R2_MC1_n180), .B(R2_MC1_n182), .Z(R2_U16_DATA2_47)
         );
  XOR2_X1 R2_MC1_U218 ( .A(R2_n1169), .B(R2_n1161), .Z(R2_MC1_n157) );
  XOR2_X1 R2_MC1_U217 ( .A(R2_n1185), .B(R2_MC1_n157), .Z(R2_MC1_n181) );
  XOR2_X1 R2_MC1_U216 ( .A(R2_MC1_n180), .B(R2_MC1_n181), .Z(R2_U16_DATA2_48)
         );
  XOR2_X1 R2_MC1_U215 ( .A(R2_n1170), .B(R2_MC1_n147), .Z(R2_MC1_n177) );
  XOR2_X1 R2_MC1_U214 ( .A(R2_n1185), .B(R2_n1192), .Z(R2_MC1_n154) );
  XOR2_X1 R2_MC1_U213 ( .A(R2_MC1_n154), .B(R2_MC1_n179), .Z(R2_MC1_n178) );
  XOR2_X1 R2_MC1_U212 ( .A(R2_MC1_n177), .B(R2_MC1_n178), .Z(R2_U16_DATA2_49)
         );
  XOR2_X1 R2_MC1_U211 ( .A(R2_n1157), .B(R2_MC1_n176), .Z(R2_MC1_n172) );
  XOR2_X1 R2_MC1_U210 ( .A(R2_MC1_n174), .B(R2_MC1_n175), .Z(R2_MC1_n173) );
  XOR2_X1 R2_MC1_U209 ( .A(R2_MC1_n172), .B(R2_MC1_n173), .Z(R2_U16_DATA2_4)
         );
  XOR2_X1 R2_MC1_U208 ( .A(R2_n1186), .B(R2_n1178), .Z(R2_MC1_n170) );
  XOR2_X1 R2_MC1_U207 ( .A(R2_n1171), .B(R2_n1163), .Z(R2_MC1_n149) );
  XOR2_X1 R2_MC1_U206 ( .A(R2_n1187), .B(R2_MC1_n149), .Z(R2_MC1_n171) );
  XOR2_X1 R2_MC1_U205 ( .A(R2_MC1_n170), .B(R2_MC1_n171), .Z(R2_U16_DATA2_50)
         );
  XOR2_X1 R2_MC1_U204 ( .A(R2_n1187), .B(R2_n1192), .Z(R2_MC1_n144) );
  XOR2_X1 R2_MC1_U203 ( .A(R2_MC1_n167), .B(R2_MC1_n168), .Z(R2_U16_DATA2_51)
         );
  XOR2_X1 R2_MC1_U202 ( .A(R2_n1173), .B(R2_MC1_n134), .Z(R2_MC1_n164) );
  XOR2_X1 R2_MC1_U201 ( .A(R2_n1188), .B(R2_n1192), .Z(R2_MC1_n139) );
  XOR2_X1 R2_MC1_U200 ( .A(R2_MC1_n139), .B(R2_MC1_n166), .Z(R2_MC1_n165) );
  XOR2_X1 R2_MC1_U199 ( .A(R2_MC1_n164), .B(R2_MC1_n165), .Z(R2_U16_DATA2_52)
         );
  XOR2_X1 R2_MC1_U198 ( .A(R2_n1189), .B(R2_n1181), .Z(R2_MC1_n162) );
  XOR2_X1 R2_MC1_U197 ( .A(R2_n1174), .B(R2_MC1_n131), .Z(R2_MC1_n163) );
  XOR2_X1 R2_MC1_U196 ( .A(R2_MC1_n162), .B(R2_MC1_n163), .Z(R2_U16_DATA2_53)
         );
  XOR2_X1 R2_MC1_U195 ( .A(R2_n1190), .B(R2_n1182), .Z(R2_MC1_n160) );
  XOR2_X1 R2_MC1_U194 ( .A(R2_n1175), .B(R2_MC1_n128), .Z(R2_MC1_n161) );
  XOR2_X1 R2_MC1_U193 ( .A(R2_MC1_n160), .B(R2_MC1_n161), .Z(R2_U16_DATA2_54)
         );
  XOR2_X1 R2_MC1_U192 ( .A(R2_n1192), .B(R2_n1191), .Z(R2_MC1_n158) );
  XOR2_X1 R2_MC1_U191 ( .A(R2_n1183), .B(R2_MC1_n126), .Z(R2_MC1_n159) );
  XOR2_X1 R2_MC1_U190 ( .A(R2_MC1_n158), .B(R2_MC1_n159), .Z(R2_U16_DATA2_55)
         );
  XOR2_X1 R2_MC1_U189 ( .A(R2_n1192), .B(R2_n1168), .Z(R2_MC1_n155) );
  XOR2_X1 R2_MC1_U188 ( .A(R2_n1177), .B(R2_MC1_n157), .Z(R2_MC1_n156) );
  XOR2_X1 R2_MC1_U187 ( .A(R2_MC1_n155), .B(R2_MC1_n156), .Z(R2_U16_DATA2_56)
         );
  XOR2_X1 R2_MC1_U186 ( .A(R2_n1162), .B(R2_MC1_n154), .Z(R2_MC1_n150) );
  XOR2_X1 R2_MC1_U185 ( .A(R2_MC1_n152), .B(R2_MC1_n153), .Z(R2_MC1_n151) );
  XOR2_X1 R2_MC1_U184 ( .A(R2_MC1_n150), .B(R2_MC1_n151), .Z(R2_U16_DATA2_57)
         );
  XOR2_X1 R2_MC1_U183 ( .A(R2_n1179), .B(R2_MC1_n149), .Z(R2_MC1_n148) );
  XOR2_X1 R2_MC1_U182 ( .A(R2_MC1_n147), .B(R2_MC1_n148), .Z(R2_U16_DATA2_58)
         );
  XOR2_X1 R2_MC1_U180 ( .A(R2_MC1_n11), .B(R2_MC1_n143), .Z(R2_U16_DATA2_59)
         );
  XOR2_X1 R2_MC1_U179 ( .A(R2_n1133), .B(R2_n1158), .Z(R2_MC1_n140) );
  XOR2_X1 R2_MC1_U178 ( .A(R2_n1141), .B(R2_MC1_n142), .Z(R2_MC1_n141) );
  XOR2_X1 R2_MC1_U177 ( .A(R2_MC1_n140), .B(R2_MC1_n141), .Z(R2_U16_DATA2_5)
         );
  XOR2_X1 R2_MC1_U176 ( .A(R2_n1165), .B(R2_MC1_n139), .Z(R2_MC1_n135) );
  XOR2_X1 R2_MC1_U175 ( .A(R2_MC1_n137), .B(R2_MC1_n138), .Z(R2_MC1_n136) );
  XOR2_X1 R2_MC1_U174 ( .A(R2_MC1_n135), .B(R2_MC1_n136), .Z(R2_U16_DATA2_60)
         );
  XOR2_X1 R2_MC1_U173 ( .A(R2_n1166), .B(R2_MC1_n134), .Z(R2_MC1_n133) );
  XOR2_X1 R2_MC1_U172 ( .A(R2_MC1_n132), .B(R2_MC1_n133), .Z(R2_U16_DATA2_61)
         );
  XOR2_X1 R2_MC1_U171 ( .A(R2_n1167), .B(R2_MC1_n131), .Z(R2_MC1_n130) );
  XOR2_X1 R2_MC1_U170 ( .A(R2_MC1_n129), .B(R2_MC1_n130), .Z(R2_U16_DATA2_62)
         );
  XOR2_X1 R2_MC1_U169 ( .A(R2_n1184), .B(R2_MC1_n128), .Z(R2_MC1_n127) );
  XOR2_X1 R2_MC1_U168 ( .A(R2_MC1_n126), .B(R2_MC1_n127), .Z(R2_U16_DATA2_63)
         );
  XOR2_X1 R2_MC1_U167 ( .A(R2_n1217), .B(R2_n1209), .Z(R2_MC1_n106) );
  XOR2_X1 R2_MC1_U166 ( .A(R2_n1200), .B(R2_n1208), .Z(R2_MC1_n36) );
  XOR2_X1 R2_MC1_U165 ( .A(R2_n1201), .B(R2_MC1_n36), .Z(R2_MC1_n125) );
  XOR2_X1 R2_MC1_U164 ( .A(R2_MC1_n106), .B(R2_MC1_n125), .Z(R2_U16_DATA2_64)
         );
  XOR2_X1 R2_MC1_U163 ( .A(R2_n1202), .B(R2_n1210), .Z(R2_MC1_n62) );
  XOR2_X1 R2_MC1_U162 ( .A(R2_n1218), .B(R2_MC1_n62), .Z(R2_MC1_n123) );
  XOR2_X1 R2_MC1_U161 ( .A(R2_n1193), .B(R2_n1200), .Z(R2_MC1_n63) );
  XOR2_X1 R2_MC1_U160 ( .A(R2_n1201), .B(R2_n1208), .Z(R2_MC1_n103) );
  XOR2_X1 R2_MC1_U159 ( .A(R2_MC1_n63), .B(R2_MC1_n103), .Z(R2_MC1_n124) );
  XOR2_X1 R2_MC1_U158 ( .A(R2_MC1_n123), .B(R2_MC1_n124), .Z(R2_U16_DATA2_65)
         );
  XOR2_X1 R2_MC1_U157 ( .A(R2_n1202), .B(R2_n1194), .Z(R2_MC1_n121) );
  XOR2_X1 R2_MC1_U156 ( .A(R2_n1219), .B(R2_n1211), .Z(R2_MC1_n99) );
  XOR2_X1 R2_MC1_U155 ( .A(R2_n1203), .B(R2_MC1_n99), .Z(R2_MC1_n122) );
  XOR2_X1 R2_MC1_U154 ( .A(R2_MC1_n121), .B(R2_MC1_n122), .Z(R2_U16_DATA2_66)
         );
  XOR2_X1 R2_MC1_U153 ( .A(R2_n1212), .B(R2_n1220), .Z(R2_MC1_n118) );
  XOR2_X1 R2_MC1_U152 ( .A(R2_n1200), .B(R2_n1195), .Z(R2_MC1_n120) );
  XOR2_X1 R2_MC1_U150 ( .A(R2_MC1_n53), .B(R2_MC1_n96), .Z(R2_MC1_n119) );
  XOR2_X1 R2_MC1_U149 ( .A(R2_MC1_n118), .B(R2_MC1_n119), .Z(R2_U16_DATA2_67)
         );
  XOR2_X1 R2_MC1_U148 ( .A(R2_n1205), .B(R2_n1213), .Z(R2_MC1_n47) );
  XOR2_X1 R2_MC1_U147 ( .A(R2_n1221), .B(R2_MC1_n47), .Z(R2_MC1_n116) );
  XOR2_X1 R2_MC1_U146 ( .A(R2_n1196), .B(R2_n1200), .Z(R2_MC1_n48) );
  XOR2_X1 R2_MC1_U145 ( .A(R2_n1204), .B(R2_n1208), .Z(R2_MC1_n95) );
  XOR2_X1 R2_MC1_U144 ( .A(R2_MC1_n48), .B(R2_MC1_n95), .Z(R2_MC1_n117) );
  XOR2_X1 R2_MC1_U143 ( .A(R2_MC1_n116), .B(R2_MC1_n117), .Z(R2_U16_DATA2_68)
         );
  XOR2_X1 R2_MC1_U142 ( .A(R2_n1222), .B(R2_n1205), .Z(R2_MC1_n114) );
  XOR2_X1 R2_MC1_U141 ( .A(R2_n1206), .B(R2_n1214), .Z(R2_MC1_n42) );
  XOR2_X1 R2_MC1_U140 ( .A(R2_n1197), .B(R2_MC1_n42), .Z(R2_MC1_n115) );
  XOR2_X1 R2_MC1_U139 ( .A(R2_MC1_n114), .B(R2_MC1_n115), .Z(R2_U16_DATA2_69)
         );
  XOR2_X1 R2_MC1_U138 ( .A(R2_n1134), .B(R2_n1159), .Z(R2_MC1_n111) );
  XOR2_X1 R2_MC1_U137 ( .A(R2_n1142), .B(R2_MC1_n113), .Z(R2_MC1_n112) );
  XOR2_X1 R2_MC1_U136 ( .A(R2_MC1_n111), .B(R2_MC1_n112), .Z(R2_U16_DATA2_6)
         );
  XOR2_X1 R2_MC1_U135 ( .A(R2_n1223), .B(R2_n1206), .Z(R2_MC1_n109) );
  XOR2_X1 R2_MC1_U134 ( .A(R2_n1207), .B(R2_n1215), .Z(R2_MC1_n39) );
  XOR2_X1 R2_MC1_U133 ( .A(R2_n1198), .B(R2_MC1_n39), .Z(R2_MC1_n110) );
  XOR2_X1 R2_MC1_U132 ( .A(R2_MC1_n109), .B(R2_MC1_n110), .Z(R2_U16_DATA2_70)
         );
  XOR2_X1 R2_MC1_U131 ( .A(R2_n1208), .B(R2_n1207), .Z(R2_MC1_n107) );
  XOR2_X1 R2_MC1_U130 ( .A(R2_n1216), .B(R2_n1224), .Z(R2_MC1_n85) );
  XOR2_X1 R2_MC1_U129 ( .A(R2_n1199), .B(R2_MC1_n85), .Z(R2_MC1_n108) );
  XOR2_X1 R2_MC1_U128 ( .A(R2_MC1_n107), .B(R2_MC1_n108), .Z(R2_U16_DATA2_71)
         );
  XOR2_X1 R2_MC1_U127 ( .A(R2_n1216), .B(R2_n1208), .Z(R2_MC1_n104) );
  XOR2_X1 R2_MC1_U126 ( .A(R2_n1193), .B(R2_MC1_n106), .Z(R2_MC1_n105) );
  XOR2_X1 R2_MC1_U125 ( .A(R2_MC1_n104), .B(R2_MC1_n105), .Z(R2_U16_DATA2_72)
         );
  XOR2_X1 R2_MC1_U124 ( .A(R2_n1194), .B(R2_n1218), .Z(R2_MC1_n54) );
  XOR2_X1 R2_MC1_U123 ( .A(R2_n1210), .B(R2_MC1_n54), .Z(R2_MC1_n101) );
  XOR2_X1 R2_MC1_U122 ( .A(R2_n1209), .B(R2_n1216), .Z(R2_MC1_n84) );
  XOR2_X1 R2_MC1_U121 ( .A(R2_MC1_n84), .B(R2_MC1_n103), .Z(R2_MC1_n102) );
  XOR2_X1 R2_MC1_U120 ( .A(R2_MC1_n101), .B(R2_MC1_n102), .Z(R2_U16_DATA2_73)
         );
  XOR2_X1 R2_MC1_U119 ( .A(R2_n1195), .B(R2_MC1_n62), .Z(R2_MC1_n100) );
  XOR2_X1 R2_MC1_U118 ( .A(R2_MC1_n99), .B(R2_MC1_n100), .Z(R2_U16_DATA2_74)
         );
  XOR2_X1 R2_MC1_U117 ( .A(R2_n1216), .B(R2_n1211), .Z(R2_MC1_n98) );
  XOR2_X1 R2_MC1_U116 ( .A(R2_n1220), .B(R2_MC1_n98), .Z(R2_MC1_n79) );
  XOR2_X1 R2_MC1_U115 ( .A(R2_MC1_n52), .B(R2_MC1_n79), .Z(R2_MC1_n97) );
  XOR2_X1 R2_MC1_U114 ( .A(R2_MC1_n96), .B(R2_MC1_n97), .Z(R2_U16_DATA2_75) );
  XOR2_X1 R2_MC1_U113 ( .A(R2_n1197), .B(R2_n1221), .Z(R2_MC1_n44) );
  XOR2_X1 R2_MC1_U112 ( .A(R2_n1213), .B(R2_MC1_n44), .Z(R2_MC1_n93) );
  XOR2_X1 R2_MC1_U111 ( .A(R2_MC1_n76), .B(R2_MC1_n95), .Z(R2_MC1_n94) );
  XOR2_X1 R2_MC1_U110 ( .A(R2_MC1_n93), .B(R2_MC1_n94), .Z(R2_U16_DATA2_76) );
  XOR2_X1 R2_MC1_U109 ( .A(R2_n1198), .B(R2_n1222), .Z(R2_MC1_n41) );
  XOR2_X1 R2_MC1_U108 ( .A(R2_n1214), .B(R2_MC1_n41), .Z(R2_MC1_n92) );
  XOR2_X1 R2_MC1_U107 ( .A(R2_MC1_n47), .B(R2_MC1_n92), .Z(R2_U16_DATA2_77) );
  XOR2_X1 R2_MC1_U106 ( .A(R2_n1199), .B(R2_n1223), .Z(R2_MC1_n38) );
  XOR2_X1 R2_MC1_U105 ( .A(R2_n1215), .B(R2_MC1_n38), .Z(R2_MC1_n91) );
  XOR2_X1 R2_MC1_U104 ( .A(R2_MC1_n42), .B(R2_MC1_n91), .Z(R2_U16_DATA2_78) );
  XOR2_X1 R2_MC1_U103 ( .A(R2_n1200), .B(R2_MC1_n39), .Z(R2_MC1_n90) );
  XOR2_X1 R2_MC1_U102 ( .A(R2_MC1_n85), .B(R2_MC1_n90), .Z(R2_U16_DATA2_79) );
  XOR2_X1 R2_MC1_U101 ( .A(R2_n1135), .B(R2_n1144), .Z(R2_MC1_n87) );
  XOR2_X1 R2_MC1_U100 ( .A(R2_n1143), .B(R2_MC1_n89), .Z(R2_MC1_n88) );
  XOR2_X1 R2_MC1_U99 ( .A(R2_MC1_n87), .B(R2_MC1_n88), .Z(R2_U16_DATA2_7) );
  XOR2_X1 R2_MC1_U98 ( .A(R2_n1201), .B(R2_n1193), .Z(R2_MC1_n67) );
  XOR2_X1 R2_MC1_U97 ( .A(R2_n1217), .B(R2_MC1_n67), .Z(R2_MC1_n86) );
  XOR2_X1 R2_MC1_U96 ( .A(R2_MC1_n85), .B(R2_MC1_n86), .Z(R2_U16_DATA2_80) );
  XOR2_X1 R2_MC1_U95 ( .A(R2_n1202), .B(R2_MC1_n54), .Z(R2_MC1_n82) );
  XOR2_X1 R2_MC1_U94 ( .A(R2_n1217), .B(R2_n1224), .Z(R2_MC1_n64) );
  XOR2_X1 R2_MC1_U93 ( .A(R2_MC1_n64), .B(R2_MC1_n84), .Z(R2_MC1_n83) );
  XOR2_X1 R2_MC1_U92 ( .A(R2_MC1_n82), .B(R2_MC1_n83), .Z(R2_U16_DATA2_81) );
  XOR2_X1 R2_MC1_U91 ( .A(R2_n1218), .B(R2_n1210), .Z(R2_MC1_n80) );
  XOR2_X1 R2_MC1_U90 ( .A(R2_n1203), .B(R2_n1195), .Z(R2_MC1_n56) );
  XOR2_X1 R2_MC1_U89 ( .A(R2_n1219), .B(R2_MC1_n56), .Z(R2_MC1_n81) );
  XOR2_X1 R2_MC1_U88 ( .A(R2_MC1_n80), .B(R2_MC1_n81), .Z(R2_U16_DATA2_82) );
  XOR2_X1 R2_MC1_U87 ( .A(R2_n1219), .B(R2_n1224), .Z(R2_MC1_n51) );
  XOR2_X1 R2_MC1_U86 ( .A(R2_MC1_n77), .B(R2_MC1_n78), .Z(R2_U16_DATA2_83) );
  XOR2_X1 R2_MC1_U85 ( .A(R2_n1205), .B(R2_MC1_n44), .Z(R2_MC1_n74) );
  XOR2_X1 R2_MC1_U84 ( .A(R2_n1220), .B(R2_n1224), .Z(R2_MC1_n49) );
  XOR2_X1 R2_MC1_U83 ( .A(R2_MC1_n49), .B(R2_MC1_n76), .Z(R2_MC1_n75) );
  XOR2_X1 R2_MC1_U82 ( .A(R2_MC1_n74), .B(R2_MC1_n75), .Z(R2_U16_DATA2_84) );
  XOR2_X1 R2_MC1_U81 ( .A(R2_n1221), .B(R2_n1213), .Z(R2_MC1_n72) );
  XOR2_X1 R2_MC1_U80 ( .A(R2_n1206), .B(R2_MC1_n41), .Z(R2_MC1_n73) );
  XOR2_X1 R2_MC1_U79 ( .A(R2_MC1_n72), .B(R2_MC1_n73), .Z(R2_U16_DATA2_85) );
  XOR2_X1 R2_MC1_U78 ( .A(R2_n1222), .B(R2_n1214), .Z(R2_MC1_n70) );
  XOR2_X1 R2_MC1_U77 ( .A(R2_n1207), .B(R2_MC1_n38), .Z(R2_MC1_n71) );
  XOR2_X1 R2_MC1_U76 ( .A(R2_MC1_n70), .B(R2_MC1_n71), .Z(R2_U16_DATA2_86) );
  XOR2_X1 R2_MC1_U75 ( .A(R2_n1224), .B(R2_n1223), .Z(R2_MC1_n68) );
  XOR2_X1 R2_MC1_U74 ( .A(R2_n1215), .B(R2_MC1_n36), .Z(R2_MC1_n69) );
  XOR2_X1 R2_MC1_U73 ( .A(R2_MC1_n68), .B(R2_MC1_n69), .Z(R2_U16_DATA2_87) );
  XOR2_X1 R2_MC1_U72 ( .A(R2_n1224), .B(R2_n1200), .Z(R2_MC1_n65) );
  XOR2_X1 R2_MC1_U71 ( .A(R2_n1209), .B(R2_MC1_n67), .Z(R2_MC1_n66) );
  XOR2_X1 R2_MC1_U70 ( .A(R2_MC1_n65), .B(R2_MC1_n66), .Z(R2_U16_DATA2_88) );
  XOR2_X1 R2_MC1_U69 ( .A(R2_n1194), .B(R2_MC1_n64), .Z(R2_MC1_n60) );
  XOR2_X1 R2_MC1_U68 ( .A(R2_MC1_n62), .B(R2_MC1_n63), .Z(R2_MC1_n61) );
  XOR2_X1 R2_MC1_U67 ( .A(R2_MC1_n60), .B(R2_MC1_n61), .Z(R2_U16_DATA2_89) );
  XOR2_X1 R2_MC1_U66 ( .A(R2_n1152), .B(R2_n1144), .Z(R2_MC1_n57) );
  XOR2_X1 R2_MC1_U65 ( .A(R2_n1129), .B(R2_MC1_n59), .Z(R2_MC1_n58) );
  XOR2_X1 R2_MC1_U64 ( .A(R2_MC1_n57), .B(R2_MC1_n58), .Z(R2_U16_DATA2_8) );
  XOR2_X1 R2_MC1_U63 ( .A(R2_n1211), .B(R2_MC1_n56), .Z(R2_MC1_n55) );
  XOR2_X1 R2_MC1_U62 ( .A(R2_MC1_n54), .B(R2_MC1_n55), .Z(R2_U16_DATA2_90) );
  XOR2_X1 R2_MC1_U60 ( .A(R2_MC1_n7), .B(R2_MC1_n50), .Z(R2_U16_DATA2_91) );
  XOR2_X1 R2_MC1_U59 ( .A(R2_n1197), .B(R2_MC1_n49), .Z(R2_MC1_n45) );
  XOR2_X1 R2_MC1_U58 ( .A(R2_MC1_n47), .B(R2_MC1_n48), .Z(R2_MC1_n46) );
  XOR2_X1 R2_MC1_U57 ( .A(R2_MC1_n45), .B(R2_MC1_n46), .Z(R2_U16_DATA2_92) );
  XOR2_X1 R2_MC1_U56 ( .A(R2_n1198), .B(R2_MC1_n44), .Z(R2_MC1_n43) );
  XOR2_X1 R2_MC1_U55 ( .A(R2_MC1_n42), .B(R2_MC1_n43), .Z(R2_U16_DATA2_93) );
  XOR2_X1 R2_MC1_U54 ( .A(R2_n1199), .B(R2_MC1_n41), .Z(R2_MC1_n40) );
  XOR2_X1 R2_MC1_U53 ( .A(R2_MC1_n39), .B(R2_MC1_n40), .Z(R2_U16_DATA2_94) );
  XOR2_X1 R2_MC1_U52 ( .A(R2_n1216), .B(R2_MC1_n38), .Z(R2_MC1_n37) );
  XOR2_X1 R2_MC1_U51 ( .A(R2_MC1_n36), .B(R2_MC1_n37), .Z(R2_U16_DATA2_95) );
  XOR2_X1 R2_MC1_U50 ( .A(R2_n1233), .B(R2_MC1_n35), .Z(R2_MC1_n34) );
  XOR2_X1 R2_MC1_U49 ( .A(R2_MC1_n33), .B(R2_MC1_n34), .Z(R2_U16_DATA2_96) );
  XOR2_X1 R2_MC1_U48 ( .A(R2_n1250), .B(R2_MC1_n32), .Z(R2_MC1_n28) );
  XOR2_X1 R2_MC1_U47 ( .A(R2_MC1_n30), .B(R2_MC1_n31), .Z(R2_MC1_n29) );
  XOR2_X1 R2_MC1_U46 ( .A(R2_MC1_n28), .B(R2_MC1_n29), .Z(R2_U16_DATA2_97) );
  XOR2_X1 R2_MC1_U45 ( .A(R2_n1226), .B(R2_n1234), .Z(R2_MC1_n25) );
  XOR2_X1 R2_MC1_U44 ( .A(R2_n1235), .B(R2_MC1_n27), .Z(R2_MC1_n26) );
  XOR2_X1 R2_MC1_U43 ( .A(R2_MC1_n25), .B(R2_MC1_n26), .Z(R2_U16_DATA2_98) );
  XOR2_X1 R2_MC1_U42 ( .A(R2_n1244), .B(R2_n1252), .Z(R2_MC1_n21) );
  XOR2_X1 R2_MC1_U41 ( .A(R2_MC1_n21), .B(R2_MC1_n22), .Z(R2_U16_DATA2_99) );
  XOR2_X1 R2_MC1_U40 ( .A(R2_n1146), .B(R2_MC1_n20), .Z(R2_MC1_n16) );
  XOR2_X1 R2_MC1_U39 ( .A(R2_MC1_n18), .B(R2_MC1_n19), .Z(R2_MC1_n17) );
  XOR2_X1 R2_MC1_U38 ( .A(R2_MC1_n16), .B(R2_MC1_n17), .Z(R2_U16_DATA2_9) );
  XOR2_X1 R2_ARK1_U128 ( .A(R2_n744), .B(R2_n872), .Z(R2_n[616]) );
  XOR2_X1 R2_ARK1_U127 ( .A(R2_n844), .B(R2_n972), .Z(R2_n[716]) );
  XOR2_X1 R2_ARK1_U126 ( .A(R2_n845), .B(R2_n973), .Z(R2_n[717]) );
  XOR2_X1 R2_ARK1_U125 ( .A(R2_n846), .B(R2_n974), .Z(R2_n[718]) );
  XOR2_X1 R2_ARK1_U124 ( .A(R2_n847), .B(R2_n975), .Z(R2_n[719]) );
  XOR2_X1 R2_ARK1_U123 ( .A(R2_n848), .B(R2_n976), .Z(R2_n[720]) );
  XOR2_X1 R2_ARK1_U122 ( .A(R2_n849), .B(R2_n977), .Z(R2_n[721]) );
  XOR2_X1 R2_ARK1_U121 ( .A(R2_n850), .B(R2_n978), .Z(R2_n[722]) );
  XOR2_X1 R2_ARK1_U120 ( .A(R2_n851), .B(R2_n979), .Z(R2_n[723]) );
  XOR2_X1 R2_ARK1_U119 ( .A(R2_n852), .B(R2_n980), .Z(R2_n[724]) );
  XOR2_X1 R2_ARK1_U118 ( .A(R2_n853), .B(R2_n981), .Z(R2_n[725]) );
  XOR2_X1 R2_ARK1_U117 ( .A(R2_n754), .B(R2_n882), .Z(R2_n[626]) );
  XOR2_X1 R2_ARK1_U116 ( .A(R2_n854), .B(R2_n982), .Z(R2_n[726]) );
  XOR2_X1 R2_ARK1_U115 ( .A(R2_n855), .B(R2_n983), .Z(R2_n[727]) );
  XOR2_X1 R2_ARK1_U114 ( .A(R2_n856), .B(R2_n984), .Z(R2_n[728]) );
  XOR2_X1 R2_ARK1_U113 ( .A(R2_n857), .B(R2_n985), .Z(R2_n[729]) );
  XOR2_X1 R2_ARK1_U112 ( .A(R2_n858), .B(R2_n986), .Z(R2_n[730]) );
  XOR2_X1 R2_ARK1_U111 ( .A(R2_n859), .B(R2_n987), .Z(R2_n[731]) );
  XOR2_X1 R2_ARK1_U110 ( .A(R2_n860), .B(R2_n988), .Z(R2_n[732]) );
  XOR2_X1 R2_ARK1_U109 ( .A(R2_n861), .B(R2_n989), .Z(R2_n[733]) );
  XOR2_X1 R2_ARK1_U108 ( .A(R2_n862), .B(R2_n990), .Z(R2_n[734]) );
  XOR2_X1 R2_ARK1_U107 ( .A(R2_n863), .B(R2_n991), .Z(R2_n[735]) );
  XOR2_X1 R2_ARK1_U106 ( .A(R2_n755), .B(R2_n883), .Z(R2_n[627]) );
  XOR2_X1 R2_ARK1_U105 ( .A(R2_n864), .B(R2_n992), .Z(R2_n[736]) );
  XOR2_X1 R2_ARK1_U104 ( .A(R2_n865), .B(R2_n993), .Z(R2_n[737]) );
  XOR2_X1 R2_ARK1_U103 ( .A(R2_n866), .B(R2_n994), .Z(R2_n[738]) );
  XOR2_X1 R2_ARK1_U102 ( .A(R2_n867), .B(R2_n995), .Z(R2_n[739]) );
  XOR2_X1 R2_ARK1_U101 ( .A(R2_n868), .B(R2_n996), .Z(R2_n[740]) );
  XOR2_X1 R2_ARK1_U100 ( .A(R2_n869), .B(R2_n997), .Z(R2_n[741]) );
  XOR2_X1 R2_ARK1_U99 ( .A(R2_n870), .B(R2_n998), .Z(R2_n[742]) );
  XOR2_X1 R2_ARK1_U98 ( .A(R2_n871), .B(R2_n999), .Z(R2_n[743]) );
  XOR2_X1 R2_ARK1_U97 ( .A(R2_n756), .B(R2_n884), .Z(R2_n[628]) );
  XOR2_X1 R2_ARK1_U96 ( .A(R2_n757), .B(R2_n885), .Z(R2_n[629]) );
  XOR2_X1 R2_ARK1_U95 ( .A(R2_n758), .B(R2_n886), .Z(R2_n[630]) );
  XOR2_X1 R2_ARK1_U94 ( .A(R2_n759), .B(R2_n887), .Z(R2_n[631]) );
  XOR2_X1 R2_ARK1_U93 ( .A(R2_n760), .B(R2_n888), .Z(R2_n[632]) );
  XOR2_X1 R2_ARK1_U92 ( .A(R2_n761), .B(R2_n889), .Z(R2_n[633]) );
  XOR2_X1 R2_ARK1_U91 ( .A(R2_n762), .B(R2_n890), .Z(R2_n[634]) );
  XOR2_X1 R2_ARK1_U90 ( .A(R2_n763), .B(R2_n891), .Z(R2_n[635]) );
  XOR2_X1 R2_ARK1_U89 ( .A(R2_n745), .B(R2_n873), .Z(R2_n[617]) );
  XOR2_X1 R2_ARK1_U88 ( .A(R2_n764), .B(R2_n892), .Z(R2_n[636]) );
  XOR2_X1 R2_ARK1_U87 ( .A(R2_n765), .B(R2_n893), .Z(R2_n[637]) );
  XOR2_X1 R2_ARK1_U86 ( .A(R2_n766), .B(R2_n894), .Z(R2_n[638]) );
  XOR2_X1 R2_ARK1_U85 ( .A(R2_n767), .B(R2_n895), .Z(R2_n[639]) );
  XOR2_X1 R2_ARK1_U84 ( .A(R2_n768), .B(R2_n896), .Z(R2_n[640]) );
  XOR2_X1 R2_ARK1_U83 ( .A(R2_n769), .B(R2_n897), .Z(R2_n[641]) );
  XOR2_X1 R2_ARK1_U82 ( .A(R2_n770), .B(R2_n898), .Z(R2_n[642]) );
  XOR2_X1 R2_ARK1_U81 ( .A(R2_n771), .B(R2_n899), .Z(R2_n[643]) );
  XOR2_X1 R2_ARK1_U80 ( .A(R2_n772), .B(R2_n900), .Z(R2_n[644]) );
  XOR2_X1 R2_ARK1_U79 ( .A(R2_n773), .B(R2_n901), .Z(R2_n[645]) );
  XOR2_X1 R2_ARK1_U78 ( .A(R2_n746), .B(R2_n874), .Z(R2_n[618]) );
  XOR2_X1 R2_ARK1_U77 ( .A(R2_n774), .B(R2_n902), .Z(R2_n[646]) );
  XOR2_X1 R2_ARK1_U76 ( .A(R2_n775), .B(R2_n903), .Z(R2_n[647]) );
  XOR2_X1 R2_ARK1_U75 ( .A(R2_n776), .B(R2_n904), .Z(R2_n[648]) );
  XOR2_X1 R2_ARK1_U74 ( .A(R2_n777), .B(R2_n905), .Z(R2_n[649]) );
  XOR2_X1 R2_ARK1_U73 ( .A(R2_n778), .B(R2_n906), .Z(R2_n[650]) );
  XOR2_X1 R2_ARK1_U72 ( .A(R2_n779), .B(R2_n907), .Z(R2_n[651]) );
  XOR2_X1 R2_ARK1_U71 ( .A(R2_n780), .B(R2_n908), .Z(R2_n[652]) );
  XOR2_X1 R2_ARK1_U70 ( .A(R2_n781), .B(R2_n909), .Z(R2_n[653]) );
  XOR2_X1 R2_ARK1_U69 ( .A(R2_n782), .B(R2_n910), .Z(R2_n[654]) );
  XOR2_X1 R2_ARK1_U68 ( .A(R2_n783), .B(R2_n911), .Z(R2_n[655]) );
  XOR2_X1 R2_ARK1_U67 ( .A(R2_n747), .B(R2_n875), .Z(R2_n[619]) );
  XOR2_X1 R2_ARK1_U66 ( .A(R2_n784), .B(R2_n912), .Z(R2_n[656]) );
  XOR2_X1 R2_ARK1_U65 ( .A(R2_n785), .B(R2_n913), .Z(R2_n[657]) );
  XOR2_X1 R2_ARK1_U64 ( .A(R2_n786), .B(R2_n914), .Z(R2_n[658]) );
  XOR2_X1 R2_ARK1_U63 ( .A(R2_n787), .B(R2_n915), .Z(R2_n[659]) );
  XOR2_X1 R2_ARK1_U62 ( .A(R2_n788), .B(R2_n916), .Z(R2_n[660]) );
  XOR2_X1 R2_ARK1_U61 ( .A(R2_n789), .B(R2_n917), .Z(R2_n[661]) );
  XOR2_X1 R2_ARK1_U60 ( .A(R2_n790), .B(R2_n918), .Z(R2_n[662]) );
  XOR2_X1 R2_ARK1_U59 ( .A(R2_n791), .B(R2_n919), .Z(R2_n[663]) );
  XOR2_X1 R2_ARK1_U58 ( .A(R2_n792), .B(R2_n920), .Z(R2_n[664]) );
  XOR2_X1 R2_ARK1_U57 ( .A(R2_n793), .B(R2_n921), .Z(R2_n[665]) );
  XOR2_X1 R2_ARK1_U56 ( .A(R2_n748), .B(R2_n876), .Z(R2_n[620]) );
  XOR2_X1 R2_ARK1_U55 ( .A(R2_n794), .B(R2_n922), .Z(R2_n[666]) );
  XOR2_X1 R2_ARK1_U54 ( .A(R2_n795), .B(R2_n923), .Z(R2_n[667]) );
  XOR2_X1 R2_ARK1_U53 ( .A(R2_n796), .B(R2_n924), .Z(R2_n[668]) );
  XOR2_X1 R2_ARK1_U52 ( .A(R2_n797), .B(R2_n925), .Z(R2_n[669]) );
  XOR2_X1 R2_ARK1_U51 ( .A(R2_n798), .B(R2_n926), .Z(R2_n[670]) );
  XOR2_X1 R2_ARK1_U50 ( .A(R2_n799), .B(R2_n927), .Z(R2_n[671]) );
  XOR2_X1 R2_ARK1_U49 ( .A(R2_n800), .B(R2_n928), .Z(R2_n[672]) );
  XOR2_X1 R2_ARK1_U48 ( .A(R2_n801), .B(R2_n929), .Z(R2_n[673]) );
  XOR2_X1 R2_ARK1_U47 ( .A(R2_n802), .B(R2_n930), .Z(R2_n[674]) );
  XOR2_X1 R2_ARK1_U46 ( .A(R2_n803), .B(R2_n931), .Z(R2_n[675]) );
  XOR2_X1 R2_ARK1_U45 ( .A(R2_n749), .B(R2_n877), .Z(R2_n[621]) );
  XOR2_X1 R2_ARK1_U44 ( .A(R2_n804), .B(R2_n932), .Z(R2_n[676]) );
  XOR2_X1 R2_ARK1_U43 ( .A(R2_n805), .B(R2_n933), .Z(R2_n[677]) );
  XOR2_X1 R2_ARK1_U42 ( .A(R2_n806), .B(R2_n934), .Z(R2_n[678]) );
  XOR2_X1 R2_ARK1_U41 ( .A(R2_n807), .B(R2_n935), .Z(R2_n[679]) );
  XOR2_X1 R2_ARK1_U40 ( .A(R2_n808), .B(R2_n936), .Z(R2_n[680]) );
  XOR2_X1 R2_ARK1_U39 ( .A(R2_n809), .B(R2_n937), .Z(R2_n[681]) );
  XOR2_X1 R2_ARK1_U38 ( .A(R2_n810), .B(R2_n938), .Z(R2_n[682]) );
  XOR2_X1 R2_ARK1_U37 ( .A(R2_n811), .B(R2_n939), .Z(R2_n[683]) );
  XOR2_X1 R2_ARK1_U36 ( .A(R2_n812), .B(R2_n940), .Z(R2_n[684]) );
  XOR2_X1 R2_ARK1_U35 ( .A(R2_n813), .B(R2_n941), .Z(R2_n[685]) );
  XOR2_X1 R2_ARK1_U34 ( .A(R2_n750), .B(R2_n878), .Z(R2_n[622]) );
  XOR2_X1 R2_ARK1_U33 ( .A(R2_n814), .B(R2_n942), .Z(R2_n[686]) );
  XOR2_X1 R2_ARK1_U32 ( .A(R2_n815), .B(R2_n943), .Z(R2_n[687]) );
  XOR2_X1 R2_ARK1_U31 ( .A(R2_n816), .B(R2_n944), .Z(R2_n[688]) );
  XOR2_X1 R2_ARK1_U30 ( .A(R2_n817), .B(R2_n945), .Z(R2_n[689]) );
  XOR2_X1 R2_ARK1_U29 ( .A(R2_n818), .B(R2_n946), .Z(R2_n[690]) );
  XOR2_X1 R2_ARK1_U28 ( .A(R2_n819), .B(R2_n947), .Z(R2_n[691]) );
  XOR2_X1 R2_ARK1_U27 ( .A(R2_n820), .B(R2_n948), .Z(R2_n[692]) );
  XOR2_X1 R2_ARK1_U26 ( .A(R2_n821), .B(R2_n949), .Z(R2_n[693]) );
  XOR2_X1 R2_ARK1_U25 ( .A(R2_n822), .B(R2_n950), .Z(R2_n[694]) );
  XOR2_X1 R2_ARK1_U24 ( .A(R2_n823), .B(R2_n951), .Z(R2_n[695]) );
  XOR2_X1 R2_ARK1_U23 ( .A(R2_n751), .B(R2_n879), .Z(R2_n[623]) );
  XOR2_X1 R2_ARK1_U22 ( .A(R2_n824), .B(R2_n952), .Z(R2_n[696]) );
  XOR2_X1 R2_ARK1_U21 ( .A(R2_n825), .B(R2_n953), .Z(R2_n[697]) );
  XOR2_X1 R2_ARK1_U20 ( .A(R2_n826), .B(R2_n954), .Z(R2_n[698]) );
  XOR2_X1 R2_ARK1_U19 ( .A(R2_n827), .B(R2_n955), .Z(R2_n[699]) );
  XOR2_X1 R2_ARK1_U18 ( .A(R2_n828), .B(R2_n956), .Z(R2_n[700]) );
  XOR2_X1 R2_ARK1_U17 ( .A(R2_n829), .B(R2_n957), .Z(R2_n[701]) );
  XOR2_X1 R2_ARK1_U16 ( .A(R2_n830), .B(R2_n958), .Z(R2_n[702]) );
  XOR2_X1 R2_ARK1_U15 ( .A(R2_n831), .B(R2_n959), .Z(R2_n[703]) );
  XOR2_X1 R2_ARK1_U14 ( .A(R2_n832), .B(R2_n960), .Z(R2_n[704]) );
  XOR2_X1 R2_ARK1_U13 ( .A(R2_n833), .B(R2_n961), .Z(R2_n[705]) );
  XOR2_X1 R2_ARK1_U12 ( .A(R2_n752), .B(R2_n880), .Z(R2_n[624]) );
  XOR2_X1 R2_ARK1_U11 ( .A(R2_n834), .B(R2_n962), .Z(R2_n[706]) );
  XOR2_X1 R2_ARK1_U10 ( .A(R2_n835), .B(R2_n963), .Z(R2_n[707]) );
  XOR2_X1 R2_ARK1_U9 ( .A(R2_n836), .B(R2_n964), .Z(R2_n[708]) );
  XOR2_X1 R2_ARK1_U8 ( .A(R2_n837), .B(R2_n965), .Z(R2_n[709]) );
  XOR2_X1 R2_ARK1_U7 ( .A(R2_n838), .B(R2_n966), .Z(R2_n[710]) );
  XOR2_X1 R2_ARK1_U6 ( .A(R2_n839), .B(R2_n967), .Z(R2_n[711]) );
  XOR2_X1 R2_ARK1_U5 ( .A(R2_n840), .B(R2_n968), .Z(R2_n[712]) );
  XOR2_X1 R2_ARK1_U4 ( .A(R2_n841), .B(R2_n969), .Z(R2_n[713]) );
  XOR2_X1 R2_ARK1_U3 ( .A(R2_n842), .B(R2_n970), .Z(R2_n[714]) );
  XOR2_X1 R2_ARK1_U2 ( .A(R2_n843), .B(R2_n971), .Z(R2_n[715]) );
  XOR2_X1 R2_ARK1_U1 ( .A(R2_n753), .B(R2_n881), .Z(R2_n[625]) );
  CLKBUF_X2 EK0_U289 ( .A(EK0_n275), .Z(EK0_n567) );
  INV_X1 EK0_U288 ( .A(EK0_n568), .ZN(EK0_n569) );
  INV_X1 EK0_U4 ( .A(EK0_U9_Z_6), .ZN(EK0_n568) );
  DFF_X2 EK0_flag_reg ( .D(EK0_n315), .CK(clk), .Q(EK0_n275) );
  NOR2_X4 EK0_U287 ( .A1(EK0_n196), .A2(EK0_n200), .ZN(EK0_n264) );
  NOR2_X4 EK0_U286 ( .A1(EK0_n200), .A2(EK0_add_99_A_1_), .ZN(EK0_n305) );
  AOI22_X1 EK0_U285 ( .A1(EK0_n195), .A2(EK0_n283), .B1(EK0_n225), .B2(
        EK0_n160), .ZN(EK0_n230) );
  AOI22_X1 EK0_U284 ( .A1(EK0_n283), .A2(EK0_n234), .B1(EK0_n198), .B2(
        EK0_n168), .ZN(EK0_n239) );
  AOI22_X1 EK0_U162 ( .A1(EK0_n283), .A2(EK0_n253), .B1(EK0_n185), .B2(
        EK0_n192), .ZN(EK0_n258) );
  AOI22_X1 EK0_U161 ( .A1(EK0_n283), .A2(EK0_n243), .B1(EK0_n197), .B2(
        EK0_n176), .ZN(EK0_n248) );
  OAI221_X1 EK0_U160 ( .B1(EK0_n251), .B2(EK0_n209), .C1(EK0_n201), .C2(
        EK0_n303), .A(EK0_n304), .ZN(EK0_U9_Z_7) );
  OAI221_X1 EK0_U159 ( .B1(EK0_n251), .B2(EK0_n211), .C1(EK0_n203), .C2(
        EK0_n303), .A(EK0_n307), .ZN(EK0_U9_Z_5) );
  INV_X1 EK0_U158 ( .A(n3259), .ZN(EK0_n202) );
  INV_X1 EK0_U157 ( .A(n3255), .ZN(EK0_n206) );
  INV_X1 EK0_U156 ( .A(n3260), .ZN(EK0_n201) );
  INV_X1 EK0_U155 ( .A(n3258), .ZN(EK0_n203) );
  INV_X1 EK0_U154 ( .A(n3244), .ZN(EK0_n209) );
  INV_X1 EK0_U153 ( .A(n3242), .ZN(EK0_n211) );
  INV_X1 EK0_U152 ( .A(n3243), .ZN(EK0_n210) );
  INV_X1 EK0_U151 ( .A(n3239), .ZN(EK0_n214) );
  INV_X1 EK0_U150 ( .A(n3256), .ZN(EK0_n205) );
  INV_X1 EK0_U149 ( .A(n3257), .ZN(EK0_n204) );
  INV_X1 EK0_U148 ( .A(n3254), .ZN(EK0_n207) );
  INV_X1 EK0_U147 ( .A(n3253), .ZN(EK0_n208) );
  INV_X1 EK0_U146 ( .A(n3240), .ZN(EK0_n213) );
  INV_X1 EK0_U145 ( .A(n3241), .ZN(EK0_n212) );
  INV_X1 EK0_U144 ( .A(n3238), .ZN(EK0_n215) );
  INV_X1 EK0_U143 ( .A(n3237), .ZN(EK0_n216) );
  INV_X1 EK0_U142 ( .A(n3127), .ZN(EK0_n220) );
  NOR2_X1 EK0_U141 ( .A1(n3125), .A2(EK0_n271), .ZN(EK0_n274) );
  INV_X1 EK0_U140 ( .A(n3126), .ZN(EK0_n221) );
  INV_X1 EK0_U139 ( .A(n3125), .ZN(EK0_n222) );
  NOR3_X1 EK0_U138 ( .A1(EK0_n221), .A2(EK0_n271), .A3(EK0_n222), .ZN(EK0_n270) );
  XNOR2_X1 EK0_U137 ( .A(EK0_n193), .B(n3163), .ZN(EK0_n269) );
  XNOR2_X1 EK0_U136 ( .A(EK0_n269), .B(EK0_n270), .ZN(EK0_n153) );
  AND2_X1 EK0_U135 ( .A1(EK0_n268), .A2(n3128), .ZN(EK0_n267) );
  XNOR2_X1 EK0_U134 ( .A(EK0_n265), .B(EK0_n266), .ZN(EK0_n154) );
  NAND2_X1 EK0_U133 ( .A1(n3127), .A2(EK0_n294), .ZN(EK0_n271) );
  NOR2_X1 EK0_U132 ( .A1(EK0_n217), .A2(n3128), .ZN(EK0_n294) );
  OAI22_X1 EK0_U131 ( .A1(EK0_n217), .A2(EK0_n276), .B1(EK0_n222), .B2(
        EK0_n297), .ZN(EK0_n295) );
  INV_X1 EK0_U130 ( .A(EK0_n289), .ZN(EK0_n218) );
  OAI22_X1 EK0_U129 ( .A1(EK0_n218), .A2(EK0_n217), .B1(n3125), .B2(EK0_n297), 
        .ZN(EK0_n298) );
  NAND2_X1 EK0_U128 ( .A1(EK0_n222), .A2(EK0_n221), .ZN(EK0_n293) );
  OAI22_X1 EK0_U127 ( .A1(EK0_n217), .A2(EK0_n292), .B1(EK0_n271), .B2(
        EK0_n293), .ZN(EK0_n290) );
  OAI21_X1 EK0_U126 ( .B1(EK0_n217), .B2(EK0_n292), .A(EK0_n302), .ZN(EK0_n300) );
  INV_X1 EK0_U125 ( .A(EK0_n276), .ZN(EK0_n219) );
  AOI22_X1 EK0_U124 ( .A1(EK0_n274), .A2(n3126), .B1(EK0_n219), .B2(EK0_n268), 
        .ZN(EK0_n273) );
  XNOR2_X1 EK0_U123 ( .A(EK0_n192), .B(n3162), .ZN(EK0_n272) );
  NOR2_X1 EK0_U122 ( .A1(n3126), .A2(EK0_n271), .ZN(EK0_n288) );
  AOI22_X1 EK0_U121 ( .A1(EK0_n288), .A2(n3125), .B1(EK0_n268), .B2(EK0_n289), 
        .ZN(EK0_n287) );
  XNOR2_X1 EK0_U120 ( .A(EK0_n191), .B(n3161), .ZN(EK0_n277) );
  NOR2_X1 EK0_U119 ( .A1(n2995), .A2(EK0_n313), .ZN(EK0_U4_Z_1) );
  NAND2_X1 EK0_U118 ( .A1(EK0_n565), .A2(EK0_n261), .ZN(EK0_n263) );
  OAI21_X1 EK0_U117 ( .B1(n2995), .B2(EK0_n261), .A(EK0_n263), .ZN(EK0_n315)
         );
  NAND2_X1 EK0_U116 ( .A1(n2996), .A2(EK0_n261), .ZN(EK0_n262) );
  OAI21_X1 EK0_U115 ( .B1(n2995), .B2(EK0_n261), .A(EK0_n262), .ZN(EK0_n314)
         );
  NAND2_X1 EK0_U114 ( .A1(EK0_U4_Z_0), .A2(EK0_n196), .ZN(EK0_n225) );
  NOR2_X1 EK0_U113 ( .A1(EK0_add_99_A_0_), .A2(n2995), .ZN(EK0_U4_Z_0) );
  NOR2_X1 EK0_U112 ( .A1(n2995), .A2(EK0_n264), .ZN(EK0_n261) );
  AOI22_X1 EK0_U111 ( .A1(EK0_n195), .A2(EK0_n282), .B1(EK0_n225), .B2(
        EK0_n159), .ZN(EK0_n229) );
  INV_X1 EK0_U110 ( .A(EK0_n229), .ZN(EK0_n17) );
  AOI22_X1 EK0_U109 ( .A1(EK0_n195), .A2(EK0_n278), .B1(EK0_n225), .B2(
        EK0_n155), .ZN(EK0_n224) );
  INV_X1 EK0_U108 ( .A(EK0_n224), .ZN(EK0_n1) );
  AOI22_X1 EK0_U107 ( .A1(EK0_n195), .A2(EK0_n280), .B1(EK0_n225), .B2(
        EK0_n157), .ZN(EK0_n227) );
  INV_X1 EK0_U106 ( .A(EK0_n227), .ZN(EK0_n9) );
  AOI22_X1 EK0_U105 ( .A1(EK0_n195), .A2(EK0_n279), .B1(EK0_n225), .B2(
        EK0_n156), .ZN(EK0_n226) );
  INV_X1 EK0_U104 ( .A(EK0_n226), .ZN(EK0_n5) );
  AOI22_X1 EK0_U103 ( .A1(EK0_n282), .A2(EK0_n234), .B1(EK0_n198), .B2(
        EK0_n167), .ZN(EK0_n238) );
  INV_X1 EK0_U102 ( .A(EK0_n238), .ZN(EK0_n18) );
  AOI22_X1 EK0_U101 ( .A1(EK0_n280), .A2(EK0_n234), .B1(EK0_n198), .B2(
        EK0_n165), .ZN(EK0_n236) );
  INV_X1 EK0_U100 ( .A(EK0_n236), .ZN(EK0_n10) );
  AOI22_X1 EK0_U99 ( .A1(EK0_n279), .A2(EK0_n234), .B1(EK0_n198), .B2(EK0_n164), .ZN(EK0_n235) );
  INV_X1 EK0_U98 ( .A(EK0_n235), .ZN(EK0_n6) );
  AOI22_X1 EK0_U97 ( .A1(EK0_n278), .A2(EK0_n234), .B1(EK0_n198), .B2(EK0_n163), .ZN(EK0_n233) );
  INV_X1 EK0_U96 ( .A(EK0_n233), .ZN(EK0_n2) );
  AOI22_X1 EK0_U95 ( .A1(EK0_n195), .A2(EK0_n281), .B1(EK0_n225), .B2(EK0_n158), .ZN(EK0_n228) );
  INV_X1 EK0_U94 ( .A(EK0_n228), .ZN(EK0_n13) );
  AOI22_X1 EK0_U93 ( .A1(EK0_n195), .A2(EK0_n285), .B1(EK0_n225), .B2(EK0_n162), .ZN(EK0_n232) );
  INV_X1 EK0_U92 ( .A(EK0_n232), .ZN(EK0_n181) );
  AOI22_X1 EK0_U91 ( .A1(EK0_n195), .A2(EK0_n284), .B1(EK0_n225), .B2(EK0_n161), .ZN(EK0_n231) );
  INV_X1 EK0_U90 ( .A(EK0_n231), .ZN(EK0_n25) );
  AOI22_X1 EK0_U89 ( .A1(EK0_n285), .A2(EK0_n234), .B1(EK0_n198), .B2(EK0_n170), .ZN(EK0_n241) );
  INV_X1 EK0_U87 ( .A(EK0_n241), .ZN(EK0_n182) );
  AOI22_X1 EK0_U85 ( .A1(EK0_n281), .A2(EK0_n234), .B1(EK0_n198), .B2(EK0_n166), .ZN(EK0_n237) );
  INV_X1 EK0_U84 ( .A(EK0_n237), .ZN(EK0_n14) );
  AOI22_X1 EK0_U83 ( .A1(EK0_n284), .A2(EK0_n234), .B1(EK0_n198), .B2(EK0_n169), .ZN(EK0_n240) );
  INV_X1 EK0_U82 ( .A(EK0_n240), .ZN(EK0_n26) );
  AOI22_X1 EK0_U81 ( .A1(EK0_n281), .A2(EK0_n253), .B1(EK0_n185), .B2(EK0_n190), .ZN(EK0_n256) );
  INV_X1 EK0_U80 ( .A(EK0_n256), .ZN(EK0_n16) );
  AOI22_X1 EK0_U79 ( .A1(EK0_n281), .A2(EK0_n243), .B1(EK0_n197), .B2(EK0_n174), .ZN(EK0_n246) );
  INV_X1 EK0_U78 ( .A(EK0_n246), .ZN(EK0_n15) );
  AOI22_X1 EK0_U77 ( .A1(EK0_n285), .A2(EK0_n253), .B1(EK0_n185), .B2(EK0_n194), .ZN(EK0_n260) );
  INV_X1 EK0_U76 ( .A(EK0_n260), .ZN(EK0_n184) );
  AOI22_X1 EK0_U75 ( .A1(EK0_n284), .A2(EK0_n253), .B1(EK0_n185), .B2(EK0_n193), .ZN(EK0_n259) );
  INV_X1 EK0_U74 ( .A(EK0_n259), .ZN(EK0_n180) );
  AOI22_X1 EK0_U73 ( .A1(EK0_n282), .A2(EK0_n253), .B1(EK0_n185), .B2(EK0_n191), .ZN(EK0_n257) );
  INV_X1 EK0_U72 ( .A(EK0_n257), .ZN(EK0_n20) );
  AOI22_X1 EK0_U71 ( .A1(EK0_n280), .A2(EK0_n253), .B1(EK0_n185), .B2(EK0_n189), .ZN(EK0_n255) );
  INV_X1 EK0_U70 ( .A(EK0_n255), .ZN(EK0_n12) );
  AOI22_X1 EK0_U69 ( .A1(EK0_n279), .A2(EK0_n253), .B1(EK0_n185), .B2(EK0_n188), .ZN(EK0_n254) );
  INV_X1 EK0_U68 ( .A(EK0_n254), .ZN(EK0_n8) );
  AOI22_X1 EK0_U67 ( .A1(EK0_n278), .A2(EK0_n253), .B1(EK0_n185), .B2(EK0_n187), .ZN(EK0_n252) );
  INV_X1 EK0_U66 ( .A(EK0_n252), .ZN(EK0_n4) );
  AOI22_X1 EK0_U65 ( .A1(EK0_n285), .A2(EK0_n243), .B1(EK0_n197), .B2(EK0_n178), .ZN(EK0_n250) );
  INV_X1 EK0_U64 ( .A(EK0_n250), .ZN(EK0_n183) );
  AOI22_X1 EK0_U63 ( .A1(EK0_n284), .A2(EK0_n243), .B1(EK0_n197), .B2(EK0_n177), .ZN(EK0_n249) );
  INV_X1 EK0_U62 ( .A(EK0_n249), .ZN(EK0_n179) );
  AOI22_X1 EK0_U61 ( .A1(EK0_n282), .A2(EK0_n243), .B1(EK0_n197), .B2(EK0_n175), .ZN(EK0_n247) );
  INV_X1 EK0_U60 ( .A(EK0_n247), .ZN(EK0_n19) );
  AOI22_X1 EK0_U59 ( .A1(EK0_n280), .A2(EK0_n243), .B1(EK0_n197), .B2(EK0_n173), .ZN(EK0_n245) );
  INV_X1 EK0_U58 ( .A(EK0_n245), .ZN(EK0_n11) );
  AOI22_X1 EK0_U57 ( .A1(EK0_n279), .A2(EK0_n243), .B1(EK0_n197), .B2(EK0_n172), .ZN(EK0_n244) );
  INV_X1 EK0_U56 ( .A(EK0_n244), .ZN(EK0_n7) );
  AOI22_X1 EK0_U55 ( .A1(EK0_n278), .A2(EK0_n243), .B1(EK0_n197), .B2(EK0_n171), .ZN(EK0_n242) );
  INV_X1 EK0_U54 ( .A(EK0_n242), .ZN(EK0_n3) );
  INV_X1 EK0_U53 ( .A(EK0_n239), .ZN(EK0_n22) );
  INV_X1 EK0_U52 ( .A(EK0_n230), .ZN(EK0_n21) );
  INV_X1 EK0_U51 ( .A(EK0_n258), .ZN(EK0_n24) );
  INV_X1 EK0_U50 ( .A(EK0_n248), .ZN(EK0_n23) );
  AOI22_X1 EK0_U49 ( .A1(n3231), .A2(EK0_n305), .B1(n3247), .B2(EK0_n264), 
        .ZN(EK0_n310) );
  OAI221_X1 EK0_U48 ( .B1(EK0_n251), .B2(EK0_n214), .C1(EK0_n206), .C2(
        EK0_n303), .A(EK0_n310), .ZN(EK0_U9_Z_2) );
  AOI22_X1 EK0_U47 ( .A1(n3230), .A2(EK0_n305), .B1(n3246), .B2(EK0_n264), 
        .ZN(EK0_n311) );
  OAI221_X1 EK0_U46 ( .B1(EK0_n251), .B2(EK0_n215), .C1(EK0_n207), .C2(
        EK0_n303), .A(EK0_n311), .ZN(EK0_U9_Z_1) );
  AOI22_X1 EK0_U45 ( .A1(n3229), .A2(EK0_n305), .B1(n3245), .B2(EK0_n264), 
        .ZN(EK0_n312) );
  OAI221_X1 EK0_U44 ( .B1(EK0_n251), .B2(EK0_n216), .C1(EK0_n208), .C2(
        EK0_n303), .A(EK0_n312), .ZN(EK0_U9_Z_0) );
  AOI22_X1 EK0_U43 ( .A1(n3235), .A2(EK0_n305), .B1(n3251), .B2(EK0_n264), 
        .ZN(EK0_n306) );
  AOI22_X1 EK0_U42 ( .A1(n3236), .A2(EK0_n305), .B1(n3252), .B2(EK0_n264), 
        .ZN(EK0_n304) );
  AOI22_X1 EK0_U41 ( .A1(n3234), .A2(EK0_n305), .B1(n3250), .B2(EK0_n264), 
        .ZN(EK0_n307) );
  AOI22_X1 EK0_U40 ( .A1(n3232), .A2(EK0_n305), .B1(n3248), .B2(EK0_n264), 
        .ZN(EK0_n309) );
  AOI22_X1 EK0_U39 ( .A1(n3233), .A2(EK0_n305), .B1(n3249), .B2(EK0_n264), 
        .ZN(EK0_n308) );
  XNOR2_X1 EK0_U38 ( .A(EK0_n203), .B(EK0_n88), .ZN(EK0_n56) );
  XNOR2_X1 EK0_U37 ( .A(EK0_n204), .B(EK0_n87), .ZN(EK0_n55) );
  XNOR2_X1 EK0_U36 ( .A(EK0_n205), .B(EK0_n86), .ZN(EK0_n54) );
  XNOR2_X1 EK0_U35 ( .A(EK0_n206), .B(EK0_n85), .ZN(EK0_n53) );
  XNOR2_X1 EK0_U34 ( .A(EK0_n207), .B(EK0_n84), .ZN(EK0_n52) );
  XNOR2_X1 EK0_U33 ( .A(EK0_n208), .B(EK0_n83), .ZN(EK0_n51) );
  XNOR2_X1 EK0_U32 ( .A(EK0_n209), .B(EK0_n74), .ZN(EK0_n42) );
  XNOR2_X1 EK0_U31 ( .A(EK0_n210), .B(EK0_n73), .ZN(EK0_n41) );
  XNOR2_X1 EK0_U30 ( .A(EK0_n211), .B(EK0_n72), .ZN(EK0_n40) );
  XNOR2_X1 EK0_U29 ( .A(EK0_n212), .B(EK0_n71), .ZN(EK0_n39) );
  XNOR2_X1 EK0_U28 ( .A(EK0_n213), .B(EK0_n70), .ZN(EK0_n38) );
  XNOR2_X1 EK0_U27 ( .A(EK0_n214), .B(EK0_n69), .ZN(EK0_n37) );
  XNOR2_X1 EK0_U26 ( .A(EK0_n215), .B(EK0_n68), .ZN(EK0_n36) );
  XNOR2_X1 EK0_U25 ( .A(EK0_n216), .B(EK0_n67), .ZN(EK0_n35) );
  XNOR2_X1 EK0_U24 ( .A(EK0_n201), .B(EK0_n90), .ZN(EK0_n58) );
  XNOR2_X1 EK0_U23 ( .A(EK0_n202), .B(EK0_n89), .ZN(EK0_n57) );
  NAND2_X1 EK0_U22 ( .A1(EK0_n276), .A2(EK0_n292), .ZN(EK0_n289) );
  INV_X1 EK0_U21 ( .A(EK0_n268), .ZN(EK0_n217) );
  BUF_X1 EK0_U20 ( .A(EK0_n564), .Z(EK0_n566) );
  BUF_X1 EK0_U19 ( .A(EK0_n564), .Z(EK0_n565) );
  INV_X1 EK0_U18 ( .A(EK0_n234), .ZN(EK0_n198) );
  INV_X1 EK0_U17 ( .A(EK0_n253), .ZN(EK0_n185) );
  INV_X1 EK0_U16 ( .A(EK0_n243), .ZN(EK0_n197) );
  INV_X1 EK0_U15 ( .A(EK0_n225), .ZN(EK0_n195) );
  INV_X1 EK0_U14 ( .A(EK0_n305), .ZN(EK0_n199) );
  INV_X1 EK0_U13 ( .A(EK0_n264), .ZN(EK0_n186) );
  AND2_X1 EK0_U12 ( .A1(EK0_n199), .A2(EK0_n251), .ZN(EK0_n313) );
  NAND2_X1 EK0_U11 ( .A1(EK0_n313), .A2(EK0_n186), .ZN(EK0_n303) );
  NOR4_X1 EK0_U10 ( .A1(1'b0), .A2(1'b0), .A3(1'b0), .A4(1'b0), .ZN(EK0_n268)
         );
  NOR2_X1 EK0_U9 ( .A1(EK0_n199), .A2(n2995), .ZN(EK0_n234) );
  NOR2_X1 EK0_U8 ( .A1(EK0_n186), .A2(n2995), .ZN(EK0_n253) );
  NOR2_X1 EK0_U7 ( .A1(EK0_n251), .A2(n2995), .ZN(EK0_n243) );
  NAND2_X2 EK0_U6 ( .A1(EK0_add_99_A_1_), .A2(EK0_n200), .ZN(EK0_n251) );
  OAI221_X1 EK0_U5 ( .B1(EK0_n251), .B2(EK0_n210), .C1(EK0_n202), .C2(EK0_n303), .A(EK0_n306), .ZN(EK0_U9_Z_6) );
  CLKBUF_X1 EK0_U3 ( .A(EK0_n275), .Z(EK0_n564) );
  DLH_X1 EK0_sbox_s2_reg_7_ ( .G(1'b1), .D(EK0_U9_Z_7), .Q(EK0_n286) );
  XOR2_X1 EK0_U282 ( .A(EK0_n164), .B(n3142), .Z(EK0_n132) );
  XOR2_X1 EK0_U281 ( .A(EK0_n132), .B(n3174), .Z(EK0_n100) );
  XOR2_X1 EK0_U280 ( .A(EK0_n165), .B(n3143), .Z(EK0_n133) );
  XOR2_X1 EK0_U279 ( .A(EK0_n133), .B(n3175), .Z(EK0_n101) );
  XOR2_X1 EK0_U278 ( .A(EK0_n166), .B(n3144), .Z(EK0_n134) );
  XOR2_X1 EK0_U277 ( .A(EK0_n134), .B(n3176), .Z(EK0_n102) );
  XOR2_X1 EK0_U276 ( .A(EK0_n167), .B(n3145), .Z(EK0_n135) );
  XOR2_X1 EK0_U275 ( .A(EK0_n135), .B(n3177), .Z(EK0_n103) );
  XOR2_X1 EK0_U274 ( .A(EK0_n168), .B(n3146), .Z(EK0_n136) );
  XOR2_X1 EK0_U273 ( .A(EK0_n136), .B(n3178), .Z(EK0_n104) );
  XOR2_X1 EK0_U272 ( .A(EK0_n169), .B(n3147), .Z(EK0_n137) );
  XOR2_X1 EK0_U271 ( .A(EK0_n137), .B(n3179), .Z(EK0_n105) );
  XOR2_X1 EK0_U270 ( .A(EK0_n170), .B(n3148), .Z(EK0_n138) );
  XOR2_X1 EK0_U269 ( .A(EK0_n138), .B(n3180), .Z(EK0_n106) );
  XOR2_X1 EK0_U268 ( .A(EK0_n171), .B(n3149), .Z(EK0_n139) );
  XOR2_X1 EK0_U267 ( .A(EK0_n139), .B(n3181), .Z(EK0_n107) );
  XOR2_X1 EK0_U266 ( .A(EK0_n172), .B(n3150), .Z(EK0_n140) );
  XOR2_X1 EK0_U265 ( .A(EK0_n140), .B(n3182), .Z(EK0_n108) );
  XOR2_X1 EK0_U264 ( .A(EK0_n173), .B(n3151), .Z(EK0_n141) );
  XOR2_X1 EK0_U263 ( .A(EK0_n141), .B(n3183), .Z(EK0_n109) );
  XOR2_X1 EK0_U262 ( .A(EK0_n174), .B(n3152), .Z(EK0_n142) );
  XOR2_X1 EK0_U261 ( .A(EK0_n142), .B(n3184), .Z(EK0_n110) );
  XOR2_X1 EK0_U260 ( .A(EK0_n175), .B(n3153), .Z(EK0_n143) );
  XOR2_X1 EK0_U259 ( .A(EK0_n143), .B(n3185), .Z(EK0_n111) );
  XOR2_X1 EK0_U258 ( .A(EK0_n176), .B(n3154), .Z(EK0_n144) );
  XOR2_X1 EK0_U257 ( .A(EK0_n144), .B(n3186), .Z(EK0_n112) );
  XOR2_X1 EK0_U256 ( .A(EK0_n177), .B(n3155), .Z(EK0_n145) );
  XOR2_X1 EK0_U255 ( .A(EK0_n145), .B(n3187), .Z(EK0_n113) );
  XOR2_X1 EK0_U254 ( .A(EK0_n178), .B(n3156), .Z(EK0_n146) );
  XOR2_X1 EK0_U253 ( .A(EK0_n146), .B(n3188), .Z(EK0_n114) );
  NAND4_X1 EK0_U252 ( .A1(n3125), .A2(n3128), .A3(EK0_n221), .A4(EK0_n220), 
        .ZN(EK0_n292) );
  NAND4_X1 EK0_U251 ( .A1(n3125), .A2(EK0_n294), .A3(EK0_n221), .A4(EK0_n220), 
        .ZN(EK0_n302) );
  XOR2_X1 EK0_U250 ( .A(EK0_n187), .B(n3157), .Z(EK0_n301) );
  XOR2_X1 EK0_U249 ( .A(EK0_n300), .B(EK0_n301), .Z(EK0_n147) );
  XOR2_X1 EK0_U248 ( .A(EK0_n147), .B(n3189), .Z(EK0_n115) );
  NAND4_X1 EK0_U247 ( .A1(n3126), .A2(n3128), .A3(EK0_n222), .A4(EK0_n220), 
        .ZN(EK0_n276) );
  NAND3_X1 EK0_U246 ( .A1(EK0_n294), .A2(EK0_n220), .A3(n3126), .ZN(EK0_n297)
         );
  XOR2_X1 EK0_U245 ( .A(EK0_n188), .B(n3158), .Z(EK0_n299) );
  XOR2_X1 EK0_U244 ( .A(EK0_n298), .B(EK0_n299), .Z(EK0_n148) );
  XOR2_X1 EK0_U243 ( .A(EK0_n148), .B(n3190), .Z(EK0_n116) );
  XOR2_X1 EK0_U242 ( .A(EK0_n189), .B(n3159), .Z(EK0_n296) );
  XOR2_X1 EK0_U241 ( .A(EK0_n295), .B(EK0_n296), .Z(EK0_n149) );
  XOR2_X1 EK0_U240 ( .A(EK0_n149), .B(n3191), .Z(EK0_n117) );
  XOR2_X1 EK0_U239 ( .A(EK0_n190), .B(n3160), .Z(EK0_n291) );
  XOR2_X1 EK0_U238 ( .A(EK0_n290), .B(EK0_n291), .Z(EK0_n150) );
  XOR2_X1 EK0_U237 ( .A(EK0_n150), .B(n3192), .Z(EK0_n118) );
  XOR2_X1 EK0_U236 ( .A(EK0_n277), .B(EK0_n287), .Z(EK0_n151) );
  XOR2_X1 EK0_U235 ( .A(EK0_n151), .B(n3193), .Z(EK0_n119) );
  XOR2_X1 EK0_U234 ( .A(EK0_n272), .B(EK0_n273), .Z(EK0_n152) );
  XOR2_X1 EK0_U233 ( .A(EK0_n152), .B(n3194), .Z(EK0_n120) );
  XOR2_X1 EK0_U232 ( .A(EK0_n153), .B(n3195), .Z(EK0_n121) );
  NAND4_X1 EK0_U231 ( .A1(EK0_n221), .A2(EK0_n220), .A3(EK0_n222), .A4(
        EK0_n267), .ZN(EK0_n265) );
  XOR2_X1 EK0_U230 ( .A(EK0_n194), .B(n3164), .Z(EK0_n266) );
  XOR2_X1 EK0_U229 ( .A(EK0_n154), .B(n3196), .Z(EK0_n122) );
  XOR2_X1 EK0_U228 ( .A(EK0_n155), .B(n3133), .Z(EK0_n123) );
  XOR2_X1 EK0_U227 ( .A(EK0_n156), .B(n3134), .Z(EK0_n124) );
  XOR2_X1 EK0_U226 ( .A(EK0_n157), .B(n3135), .Z(EK0_n125) );
  XOR2_X1 EK0_U225 ( .A(EK0_n158), .B(n3136), .Z(EK0_n126) );
  XOR2_X1 EK0_U224 ( .A(EK0_n159), .B(n3137), .Z(EK0_n127) );
  XOR2_X1 EK0_U223 ( .A(EK0_n160), .B(n3138), .Z(EK0_n128) );
  XOR2_X1 EK0_U222 ( .A(EK0_n161), .B(n3139), .Z(EK0_n129) );
  XOR2_X1 EK0_U221 ( .A(EK0_n162), .B(n3140), .Z(EK0_n130) );
  XOR2_X1 EK0_U220 ( .A(EK0_n163), .B(n3141), .Z(EK0_n131) );
  XOR2_X1 EK0_U219 ( .A(EK0_n123), .B(n3165), .Z(EK0_n91) );
  XOR2_X1 EK0_U218 ( .A(EK0_n91), .B(n3197), .Z(EK0_n59) );
  XOR2_X1 EK0_U217 ( .A(n3229), .B(EK0_n59), .Z(EK0_n27) );
  XOR2_X1 EK0_U216 ( .A(EK0_n124), .B(n3166), .Z(EK0_n92) );
  XOR2_X1 EK0_U215 ( .A(EK0_n92), .B(n3198), .Z(EK0_n60) );
  XOR2_X1 EK0_U214 ( .A(n3230), .B(EK0_n60), .Z(EK0_n28) );
  XOR2_X1 EK0_U213 ( .A(EK0_n125), .B(n3167), .Z(EK0_n93) );
  XOR2_X1 EK0_U212 ( .A(EK0_n93), .B(n3199), .Z(EK0_n61) );
  XOR2_X1 EK0_U211 ( .A(n3231), .B(EK0_n61), .Z(EK0_n29) );
  XOR2_X1 EK0_U210 ( .A(EK0_n126), .B(n3168), .Z(EK0_n94) );
  XOR2_X1 EK0_U209 ( .A(EK0_n94), .B(n3200), .Z(EK0_n62) );
  XOR2_X1 EK0_U208 ( .A(n3232), .B(EK0_n62), .Z(EK0_n30) );
  XOR2_X1 EK0_U207 ( .A(EK0_n127), .B(n3169), .Z(EK0_n95) );
  XOR2_X1 EK0_U206 ( .A(EK0_n95), .B(n3201), .Z(EK0_n63) );
  XOR2_X1 EK0_U205 ( .A(n3233), .B(EK0_n63), .Z(EK0_n31) );
  XOR2_X1 EK0_U204 ( .A(EK0_n128), .B(n3170), .Z(EK0_n96) );
  XOR2_X1 EK0_U203 ( .A(EK0_n96), .B(n3202), .Z(EK0_n64) );
  XOR2_X1 EK0_U202 ( .A(n3234), .B(EK0_n64), .Z(EK0_n32) );
  XOR2_X1 EK0_U201 ( .A(EK0_n129), .B(n3171), .Z(EK0_n97) );
  XOR2_X1 EK0_U200 ( .A(EK0_n97), .B(n3203), .Z(EK0_n65) );
  XOR2_X1 EK0_U199 ( .A(n3235), .B(EK0_n65), .Z(EK0_n33) );
  XOR2_X1 EK0_U198 ( .A(EK0_n130), .B(n3172), .Z(EK0_n98) );
  XOR2_X1 EK0_U197 ( .A(EK0_n98), .B(n3204), .Z(EK0_n66) );
  XOR2_X1 EK0_U196 ( .A(n3236), .B(EK0_n66), .Z(EK0_n34) );
  XOR2_X1 EK0_U195 ( .A(EK0_n131), .B(n3173), .Z(EK0_n99) );
  XOR2_X1 EK0_U194 ( .A(EK0_n99), .B(n3205), .Z(EK0_n67) );
  XOR2_X1 EK0_U193 ( .A(EK0_n100), .B(n3206), .Z(EK0_n68) );
  XOR2_X1 EK0_U192 ( .A(EK0_n101), .B(n3207), .Z(EK0_n69) );
  XOR2_X1 EK0_U191 ( .A(EK0_n102), .B(n3208), .Z(EK0_n70) );
  XOR2_X1 EK0_U190 ( .A(EK0_n103), .B(n3209), .Z(EK0_n71) );
  XOR2_X1 EK0_U189 ( .A(EK0_n104), .B(n3210), .Z(EK0_n72) );
  XOR2_X1 EK0_U188 ( .A(EK0_n105), .B(n3211), .Z(EK0_n73) );
  XOR2_X1 EK0_U187 ( .A(EK0_n106), .B(n3212), .Z(EK0_n74) );
  XOR2_X1 EK0_U186 ( .A(EK0_n107), .B(n3213), .Z(EK0_n75) );
  XOR2_X1 EK0_U185 ( .A(n3245), .B(EK0_n75), .Z(EK0_n43) );
  XOR2_X1 EK0_U184 ( .A(EK0_n108), .B(n3214), .Z(EK0_n76) );
  XOR2_X1 EK0_U183 ( .A(n3246), .B(EK0_n76), .Z(EK0_n44) );
  XOR2_X1 EK0_U182 ( .A(EK0_n109), .B(n3215), .Z(EK0_n77) );
  XOR2_X1 EK0_U181 ( .A(n3247), .B(EK0_n77), .Z(EK0_n45) );
  XOR2_X1 EK0_U180 ( .A(EK0_n110), .B(n3216), .Z(EK0_n78) );
  XOR2_X1 EK0_U179 ( .A(n3248), .B(EK0_n78), .Z(EK0_n46) );
  XOR2_X1 EK0_U178 ( .A(EK0_n111), .B(n3217), .Z(EK0_n79) );
  XOR2_X1 EK0_U177 ( .A(n3249), .B(EK0_n79), .Z(EK0_n47) );
  XOR2_X1 EK0_U176 ( .A(EK0_n112), .B(n3218), .Z(EK0_n80) );
  XOR2_X1 EK0_U175 ( .A(n3250), .B(EK0_n80), .Z(EK0_n48) );
  XOR2_X1 EK0_U174 ( .A(EK0_n113), .B(n3219), .Z(EK0_n81) );
  XOR2_X1 EK0_U173 ( .A(n3251), .B(EK0_n81), .Z(EK0_n49) );
  XOR2_X1 EK0_U172 ( .A(EK0_n114), .B(n3220), .Z(EK0_n82) );
  XOR2_X1 EK0_U171 ( .A(n3252), .B(EK0_n82), .Z(EK0_n50) );
  XOR2_X1 EK0_U170 ( .A(EK0_n115), .B(n3221), .Z(EK0_n83) );
  XOR2_X1 EK0_U169 ( .A(EK0_n116), .B(n3222), .Z(EK0_n84) );
  XOR2_X1 EK0_U168 ( .A(EK0_n117), .B(n3223), .Z(EK0_n85) );
  XOR2_X1 EK0_U167 ( .A(EK0_n118), .B(n3224), .Z(EK0_n86) );
  XOR2_X1 EK0_U166 ( .A(EK0_n119), .B(n3225), .Z(EK0_n87) );
  XOR2_X1 EK0_U165 ( .A(EK0_n120), .B(n3226), .Z(EK0_n88) );
  XOR2_X1 EK0_U164 ( .A(EK0_n121), .B(n3227), .Z(EK0_n89) );
  XOR2_X1 EK0_U163 ( .A(EK0_n122), .B(n3228), .Z(EK0_n90) );
  OAI221_X2 EK0_U88 ( .B1(EK0_n251), .B2(EK0_n213), .C1(EK0_n205), .C2(
        EK0_n303), .A(EK0_n309), .ZN(EK0_U9_Z_3) );
  OAI221_X2 EK0_U86 ( .B1(EK0_n251), .B2(EK0_n212), .C1(EK0_n204), .C2(
        EK0_n303), .A(EK0_n308), .ZN(EK0_U9_Z_4) );
  DLH_X1 EK0_temp_expanded_key_reg_96_ ( .G(EK0_n567), .D(EK0_n27), .Q(n[3093]) );
  DLH_X1 EK0_temp_expanded_key_reg_64_ ( .G(EK0_n567), .D(EK0_n59), .Q(n[3061]) );
  DLH_X1 EK0_temp_expanded_key_reg_32_ ( .G(EK0_n567), .D(EK0_n91), .Q(n[3029]) );
  DLH_X1 EK0_temp_expanded_key_reg_0_ ( .G(EK0_n567), .D(EK0_n123), .Q(n[2997]) );
  DFF_X1 EK0_sub_word_reg_0_ ( .D(EK0_n1), .CK(clk), .Q(EK0_n155) );
  DLH_X1 EK0_temp_expanded_key_reg_97_ ( .G(EK0_n567), .D(EK0_n28), .Q(n[3094]) );
  DLH_X1 EK0_temp_expanded_key_reg_65_ ( .G(EK0_n567), .D(EK0_n60), .Q(n[3062]) );
  DLH_X1 EK0_temp_expanded_key_reg_33_ ( .G(EK0_n565), .D(EK0_n92), .Q(n[3030]) );
  DLH_X1 EK0_temp_expanded_key_reg_1_ ( .G(EK0_n567), .D(EK0_n124), .Q(n[2998]) );
  DFF_X1 EK0_sub_word_reg_1_ ( .D(EK0_n5), .CK(clk), .Q(EK0_n156) );
  DLH_X1 EK0_temp_expanded_key_reg_98_ ( .G(EK0_n567), .D(EK0_n29), .Q(n[3095]) );
  DLH_X1 EK0_temp_expanded_key_reg_66_ ( .G(EK0_n567), .D(EK0_n61), .Q(n[3063]) );
  DLH_X1 EK0_temp_expanded_key_reg_34_ ( .G(EK0_n565), .D(EK0_n93), .Q(n[3031]) );
  DLH_X1 EK0_temp_expanded_key_reg_2_ ( .G(EK0_n567), .D(EK0_n125), .Q(n[2999]) );
  DFF_X1 EK0_sub_word_reg_2_ ( .D(EK0_n9), .CK(clk), .Q(EK0_n157) );
  DLH_X1 EK0_temp_expanded_key_reg_99_ ( .G(EK0_n567), .D(EK0_n30), .Q(n[3096]) );
  DLH_X1 EK0_temp_expanded_key_reg_67_ ( .G(EK0_n565), .D(EK0_n62), .Q(n[3064]) );
  DLH_X1 EK0_temp_expanded_key_reg_35_ ( .G(EK0_n567), .D(EK0_n94), .Q(n[3032]) );
  DLH_X1 EK0_temp_expanded_key_reg_3_ ( .G(EK0_n567), .D(EK0_n126), .Q(n[3000]) );
  DFF_X1 EK0_sub_word_reg_3_ ( .D(EK0_n13), .CK(clk), .Q(EK0_n158) );
  DLH_X1 EK0_temp_expanded_key_reg_100_ ( .G(EK0_n567), .D(EK0_n31), .Q(
        n[3097]) );
  DLH_X1 EK0_temp_expanded_key_reg_68_ ( .G(EK0_n567), .D(EK0_n63), .Q(n[3065]) );
  DLH_X1 EK0_temp_expanded_key_reg_36_ ( .G(EK0_n566), .D(EK0_n95), .Q(n[3033]) );
  DLH_X1 EK0_temp_expanded_key_reg_4_ ( .G(EK0_n567), .D(EK0_n127), .Q(n[3001]) );
  DFF_X1 EK0_sub_word_reg_4_ ( .D(EK0_n17), .CK(clk), .Q(EK0_n159) );
  DLH_X1 EK0_temp_expanded_key_reg_101_ ( .G(EK0_n567), .D(EK0_n32), .Q(
        n[3098]) );
  DLH_X1 EK0_temp_expanded_key_reg_69_ ( .G(EK0_n567), .D(EK0_n64), .Q(n[3066]) );
  DLH_X1 EK0_temp_expanded_key_reg_37_ ( .G(EK0_n565), .D(EK0_n96), .Q(n[3034]) );
  DLH_X1 EK0_temp_expanded_key_reg_5_ ( .G(EK0_n567), .D(EK0_n128), .Q(n[3002]) );
  DFF_X1 EK0_sub_word_reg_5_ ( .D(EK0_n21), .CK(clk), .Q(EK0_n160) );
  DLH_X1 EK0_temp_expanded_key_reg_102_ ( .G(EK0_n567), .D(EK0_n33), .Q(
        n[3099]) );
  DLH_X1 EK0_temp_expanded_key_reg_70_ ( .G(EK0_n566), .D(EK0_n65), .Q(n[3067]) );
  DLH_X1 EK0_temp_expanded_key_reg_38_ ( .G(EK0_n567), .D(EK0_n97), .Q(n[3035]) );
  DLH_X1 EK0_temp_expanded_key_reg_6_ ( .G(EK0_n567), .D(EK0_n129), .Q(n[3003]) );
  DFF_X1 EK0_sub_word_reg_6_ ( .D(EK0_n25), .CK(clk), .Q(EK0_n161) );
  DLH_X1 EK0_temp_expanded_key_reg_103_ ( .G(EK0_n565), .D(EK0_n34), .Q(
        n[3100]) );
  DLH_X1 EK0_temp_expanded_key_reg_71_ ( .G(EK0_n566), .D(EK0_n66), .Q(n[3068]) );
  DLH_X1 EK0_temp_expanded_key_reg_39_ ( .G(EK0_n275), .D(EK0_n98), .Q(n[3036]) );
  DLH_X1 EK0_temp_expanded_key_reg_7_ ( .G(EK0_n567), .D(EK0_n130), .Q(n[3004]) );
  DFF_X1 EK0_sub_word_reg_7_ ( .D(EK0_n181), .CK(clk), .Q(EK0_n162) );
  DLH_X1 EK0_temp_expanded_key_reg_104_ ( .G(EK0_n275), .D(EK0_n35), .Q(
        n[3101]) );
  DLH_X1 EK0_temp_expanded_key_reg_72_ ( .G(EK0_n567), .D(EK0_n67), .Q(n[3069]) );
  DLH_X1 EK0_temp_expanded_key_reg_40_ ( .G(EK0_n275), .D(EK0_n99), .Q(n[3037]) );
  DLH_X1 EK0_temp_expanded_key_reg_8_ ( .G(EK0_n567), .D(EK0_n131), .Q(n[3005]) );
  DFF_X1 EK0_sub_word_reg_8_ ( .D(EK0_n2), .CK(clk), .Q(EK0_n163) );
  DLH_X1 EK0_temp_expanded_key_reg_105_ ( .G(EK0_n564), .D(EK0_n36), .Q(
        n[3102]) );
  DLH_X1 EK0_temp_expanded_key_reg_73_ ( .G(EK0_n566), .D(EK0_n68), .Q(n[3070]) );
  DLH_X1 EK0_temp_expanded_key_reg_41_ ( .G(EK0_n275), .D(EK0_n100), .Q(
        n[3038]) );
  DLH_X1 EK0_temp_expanded_key_reg_9_ ( .G(EK0_n275), .D(EK0_n132), .Q(n[3006]) );
  DFF_X1 EK0_sub_word_reg_9_ ( .D(EK0_n6), .CK(clk), .Q(EK0_n164) );
  DLH_X1 EK0_temp_expanded_key_reg_106_ ( .G(EK0_n567), .D(EK0_n37), .Q(
        n[3103]) );
  DLH_X1 EK0_temp_expanded_key_reg_74_ ( .G(EK0_n275), .D(EK0_n69), .Q(n[3071]) );
  DLH_X1 EK0_temp_expanded_key_reg_42_ ( .G(EK0_n567), .D(EK0_n101), .Q(
        n[3039]) );
  DLH_X1 EK0_temp_expanded_key_reg_10_ ( .G(EK0_n275), .D(EK0_n133), .Q(
        n[3007]) );
  DFF_X1 EK0_sub_word_reg_10_ ( .D(EK0_n10), .CK(clk), .Q(EK0_n165) );
  DLH_X1 EK0_temp_expanded_key_reg_107_ ( .G(EK0_n275), .D(EK0_n38), .Q(
        n[3104]) );
  DLH_X1 EK0_temp_expanded_key_reg_75_ ( .G(EK0_n567), .D(EK0_n70), .Q(n[3072]) );
  DLH_X1 EK0_temp_expanded_key_reg_43_ ( .G(EK0_n275), .D(EK0_n102), .Q(
        n[3040]) );
  DLH_X1 EK0_temp_expanded_key_reg_11_ ( .G(EK0_n567), .D(EK0_n134), .Q(
        n[3008]) );
  DFF_X1 EK0_sub_word_reg_11_ ( .D(EK0_n14), .CK(clk), .Q(EK0_n166) );
  DLH_X1 EK0_temp_expanded_key_reg_108_ ( .G(EK0_n567), .D(EK0_n39), .Q(
        n[3105]) );
  DLH_X1 EK0_temp_expanded_key_reg_76_ ( .G(EK0_n275), .D(EK0_n71), .Q(n[3073]) );
  DLH_X1 EK0_temp_expanded_key_reg_44_ ( .G(EK0_n567), .D(EK0_n103), .Q(
        n[3041]) );
  DLH_X1 EK0_temp_expanded_key_reg_12_ ( .G(EK0_n275), .D(EK0_n135), .Q(
        n[3009]) );
  DFF_X1 EK0_sub_word_reg_12_ ( .D(EK0_n18), .CK(clk), .Q(EK0_n167) );
  DLH_X1 EK0_temp_expanded_key_reg_109_ ( .G(EK0_n567), .D(EK0_n40), .Q(
        n[3106]) );
  DLH_X1 EK0_temp_expanded_key_reg_77_ ( .G(EK0_n275), .D(EK0_n72), .Q(n[3074]) );
  DLH_X1 EK0_temp_expanded_key_reg_45_ ( .G(EK0_n567), .D(EK0_n104), .Q(
        n[3042]) );
  DLH_X1 EK0_temp_expanded_key_reg_13_ ( .G(EK0_n566), .D(EK0_n136), .Q(
        n[3010]) );
  DFF_X1 EK0_sub_word_reg_13_ ( .D(EK0_n22), .CK(clk), .Q(EK0_n168) );
  DLH_X1 EK0_temp_expanded_key_reg_110_ ( .G(EK0_n565), .D(EK0_n41), .Q(
        n[3107]) );
  DLH_X1 EK0_temp_expanded_key_reg_78_ ( .G(EK0_n566), .D(EK0_n73), .Q(n[3075]) );
  DLH_X1 EK0_temp_expanded_key_reg_46_ ( .G(EK0_n565), .D(EK0_n105), .Q(
        n[3043]) );
  DLH_X1 EK0_temp_expanded_key_reg_14_ ( .G(EK0_n566), .D(EK0_n137), .Q(
        n[3011]) );
  DFF_X1 EK0_sub_word_reg_14_ ( .D(EK0_n26), .CK(clk), .Q(EK0_n169) );
  DLH_X1 EK0_temp_expanded_key_reg_111_ ( .G(EK0_n565), .D(EK0_n42), .Q(
        n[3108]) );
  DLH_X1 EK0_temp_expanded_key_reg_79_ ( .G(EK0_n566), .D(EK0_n74), .Q(n[3076]) );
  DLH_X1 EK0_temp_expanded_key_reg_47_ ( .G(EK0_n565), .D(EK0_n106), .Q(
        n[3044]) );
  DLH_X1 EK0_temp_expanded_key_reg_15_ ( .G(EK0_n566), .D(EK0_n138), .Q(
        n[3012]) );
  DFF_X1 EK0_sub_word_reg_15_ ( .D(EK0_n182), .CK(clk), .Q(EK0_n170) );
  DLH_X1 EK0_temp_expanded_key_reg_112_ ( .G(EK0_n566), .D(EK0_n43), .Q(
        n[3109]) );
  DLH_X1 EK0_temp_expanded_key_reg_80_ ( .G(EK0_n566), .D(EK0_n75), .Q(n[3077]) );
  DLH_X1 EK0_temp_expanded_key_reg_48_ ( .G(EK0_n565), .D(EK0_n107), .Q(
        n[3045]) );
  DLH_X1 EK0_temp_expanded_key_reg_16_ ( .G(EK0_n566), .D(EK0_n139), .Q(
        n[3013]) );
  DFF_X1 EK0_sub_word_reg_16_ ( .D(EK0_n3), .CK(clk), .Q(EK0_n171) );
  DLH_X1 EK0_temp_expanded_key_reg_113_ ( .G(EK0_n565), .D(EK0_n44), .Q(
        n[3110]) );
  DLH_X1 EK0_temp_expanded_key_reg_81_ ( .G(EK0_n565), .D(EK0_n76), .Q(n[3078]) );
  DLH_X1 EK0_temp_expanded_key_reg_49_ ( .G(EK0_n566), .D(EK0_n108), .Q(
        n[3046]) );
  DLH_X1 EK0_temp_expanded_key_reg_17_ ( .G(EK0_n565), .D(EK0_n140), .Q(
        n[3014]) );
  DFF_X1 EK0_sub_word_reg_17_ ( .D(EK0_n7), .CK(clk), .Q(EK0_n172) );
  DLH_X1 EK0_temp_expanded_key_reg_114_ ( .G(EK0_n566), .D(EK0_n45), .Q(
        n[3111]) );
  DLH_X1 EK0_temp_expanded_key_reg_82_ ( .G(EK0_n565), .D(EK0_n77), .Q(n[3079]) );
  DLH_X1 EK0_temp_expanded_key_reg_50_ ( .G(EK0_n566), .D(EK0_n109), .Q(
        n[3047]) );
  DLH_X1 EK0_temp_expanded_key_reg_18_ ( .G(EK0_n565), .D(EK0_n141), .Q(
        n[3015]) );
  DFF_X1 EK0_sub_word_reg_18_ ( .D(EK0_n11), .CK(clk), .Q(EK0_n173) );
  DLH_X1 EK0_temp_expanded_key_reg_115_ ( .G(EK0_n566), .D(EK0_n46), .Q(
        n[3112]) );
  DLH_X1 EK0_temp_expanded_key_reg_83_ ( .G(EK0_n565), .D(EK0_n78), .Q(n[3080]) );
  DLH_X1 EK0_temp_expanded_key_reg_51_ ( .G(EK0_n566), .D(EK0_n110), .Q(
        n[3048]) );
  DLH_X1 EK0_temp_expanded_key_reg_19_ ( .G(EK0_n565), .D(EK0_n142), .Q(
        n[3016]) );
  DFF_X1 EK0_sub_word_reg_19_ ( .D(EK0_n15), .CK(clk), .Q(EK0_n174) );
  DLH_X1 EK0_temp_expanded_key_reg_116_ ( .G(EK0_n275), .D(EK0_n47), .Q(
        n[3113]) );
  DLH_X1 EK0_temp_expanded_key_reg_84_ ( .G(EK0_n275), .D(EK0_n79), .Q(n[3081]) );
  DLH_X1 EK0_temp_expanded_key_reg_52_ ( .G(EK0_n275), .D(EK0_n111), .Q(
        n[3049]) );
  DLH_X1 EK0_temp_expanded_key_reg_20_ ( .G(EK0_n275), .D(EK0_n143), .Q(
        n[3017]) );
  DFF_X1 EK0_sub_word_reg_20_ ( .D(EK0_n19), .CK(clk), .Q(EK0_n175) );
  DLH_X1 EK0_temp_expanded_key_reg_117_ ( .G(EK0_n275), .D(EK0_n48), .Q(
        n[3114]) );
  DLH_X1 EK0_temp_expanded_key_reg_85_ ( .G(EK0_n275), .D(EK0_n80), .Q(n[3082]) );
  DLH_X1 EK0_temp_expanded_key_reg_53_ ( .G(EK0_n275), .D(EK0_n112), .Q(
        n[3050]) );
  DLH_X1 EK0_temp_expanded_key_reg_21_ ( .G(EK0_n275), .D(EK0_n144), .Q(
        n[3018]) );
  DFF_X1 EK0_sub_word_reg_21_ ( .D(EK0_n23), .CK(clk), .Q(EK0_n176) );
  DLH_X1 EK0_temp_expanded_key_reg_118_ ( .G(EK0_n275), .D(EK0_n49), .Q(
        n[3115]) );
  DLH_X1 EK0_temp_expanded_key_reg_86_ ( .G(EK0_n275), .D(EK0_n81), .Q(n[3083]) );
  DLH_X1 EK0_temp_expanded_key_reg_54_ ( .G(EK0_n275), .D(EK0_n113), .Q(
        n[3051]) );
  DLH_X1 EK0_temp_expanded_key_reg_22_ ( .G(EK0_n275), .D(EK0_n145), .Q(
        n[3019]) );
  DFF_X1 EK0_sub_word_reg_22_ ( .D(EK0_n179), .CK(clk), .Q(EK0_n177) );
  DLH_X1 EK0_temp_expanded_key_reg_119_ ( .G(EK0_n564), .D(EK0_n50), .Q(
        n[3116]) );
  DLH_X1 EK0_temp_expanded_key_reg_87_ ( .G(EK0_n564), .D(EK0_n82), .Q(n[3084]) );
  DLH_X1 EK0_temp_expanded_key_reg_55_ ( .G(EK0_n564), .D(EK0_n114), .Q(
        n[3052]) );
  DLH_X1 EK0_temp_expanded_key_reg_23_ ( .G(EK0_n564), .D(EK0_n146), .Q(
        n[3020]) );
  DFF_X1 EK0_sub_word_reg_23_ ( .D(EK0_n183), .CK(clk), .Q(EK0_n178) );
  DLH_X1 EK0_temp_expanded_key_reg_120_ ( .G(EK0_n275), .D(EK0_n51), .Q(
        n[3117]) );
  DLH_X1 EK0_temp_expanded_key_reg_88_ ( .G(EK0_n275), .D(EK0_n83), .Q(n[3085]) );
  DLH_X1 EK0_temp_expanded_key_reg_56_ ( .G(EK0_n564), .D(EK0_n115), .Q(
        n[3053]) );
  DLH_X1 EK0_temp_expanded_key_reg_24_ ( .G(EK0_n564), .D(EK0_n147), .Q(
        n[3021]) );
  DFF_X1 EK0_sub_word_reg_24_ ( .D(EK0_n4), .CK(clk), .Q(EK0_n187) );
  DLH_X1 EK0_temp_expanded_key_reg_121_ ( .G(EK0_n275), .D(EK0_n52), .Q(
        n[3118]) );
  DLH_X1 EK0_temp_expanded_key_reg_89_ ( .G(EK0_n275), .D(EK0_n84), .Q(n[3086]) );
  DLH_X1 EK0_temp_expanded_key_reg_57_ ( .G(EK0_n275), .D(EK0_n116), .Q(
        n[3054]) );
  DLH_X1 EK0_temp_expanded_key_reg_25_ ( .G(EK0_n275), .D(EK0_n148), .Q(
        n[3022]) );
  DFF_X1 EK0_sub_word_reg_25_ ( .D(EK0_n8), .CK(clk), .Q(EK0_n188) );
  DLH_X1 EK0_temp_expanded_key_reg_122_ ( .G(EK0_n275), .D(EK0_n53), .Q(
        n[3119]) );
  DLH_X1 EK0_temp_expanded_key_reg_90_ ( .G(EK0_n565), .D(EK0_n85), .Q(n[3087]) );
  DLH_X1 EK0_temp_expanded_key_reg_58_ ( .G(EK0_n566), .D(EK0_n117), .Q(
        n[3055]) );
  DLH_X1 EK0_temp_expanded_key_reg_26_ ( .G(EK0_n565), .D(EK0_n149), .Q(
        n[3023]) );
  DFF_X1 EK0_sub_word_reg_26_ ( .D(EK0_n12), .CK(clk), .Q(EK0_n189) );
  DLH_X1 EK0_temp_expanded_key_reg_123_ ( .G(EK0_n566), .D(EK0_n54), .Q(
        n[3120]) );
  DLH_X1 EK0_temp_expanded_key_reg_91_ ( .G(EK0_n565), .D(EK0_n86), .Q(n[3088]) );
  DLH_X1 EK0_temp_expanded_key_reg_59_ ( .G(EK0_n566), .D(EK0_n118), .Q(
        n[3056]) );
  DLH_X1 EK0_temp_expanded_key_reg_27_ ( .G(EK0_n565), .D(EK0_n150), .Q(
        n[3024]) );
  DFF_X1 EK0_sub_word_reg_27_ ( .D(EK0_n16), .CK(clk), .Q(EK0_n190) );
  DLH_X1 EK0_temp_expanded_key_reg_124_ ( .G(EK0_n566), .D(EK0_n55), .Q(
        n[3121]) );
  DLH_X1 EK0_temp_expanded_key_reg_92_ ( .G(EK0_n566), .D(EK0_n87), .Q(n[3089]) );
  DLH_X1 EK0_temp_expanded_key_reg_60_ ( .G(EK0_n565), .D(EK0_n119), .Q(
        n[3057]) );
  DLH_X1 EK0_temp_expanded_key_reg_28_ ( .G(EK0_n566), .D(EK0_n151), .Q(
        n[3025]) );
  DFF_X1 EK0_sub_word_reg_28_ ( .D(EK0_n20), .CK(clk), .Q(EK0_n191) );
  DLH_X1 EK0_temp_expanded_key_reg_125_ ( .G(EK0_n565), .D(EK0_n56), .Q(
        n[3122]) );
  DLH_X1 EK0_temp_expanded_key_reg_93_ ( .G(EK0_n566), .D(EK0_n88), .Q(n[3090]) );
  DLH_X1 EK0_temp_expanded_key_reg_61_ ( .G(EK0_n565), .D(EK0_n120), .Q(
        n[3058]) );
  DLH_X1 EK0_temp_expanded_key_reg_29_ ( .G(EK0_n566), .D(EK0_n152), .Q(
        n[3026]) );
  DFF_X1 EK0_sub_word_reg_29_ ( .D(EK0_n24), .CK(clk), .Q(EK0_n192) );
  DLH_X1 EK0_temp_expanded_key_reg_126_ ( .G(EK0_n565), .D(EK0_n57), .Q(
        n[3123]) );
  DLH_X1 EK0_temp_expanded_key_reg_94_ ( .G(EK0_n566), .D(EK0_n89), .Q(n[3091]) );
  DLH_X1 EK0_temp_expanded_key_reg_62_ ( .G(EK0_n565), .D(EK0_n121), .Q(
        n[3059]) );
  DLH_X1 EK0_temp_expanded_key_reg_30_ ( .G(EK0_n566), .D(EK0_n153), .Q(
        n[3027]) );
  DFF_X1 EK0_sub_word_reg_30_ ( .D(EK0_n180), .CK(clk), .Q(EK0_n193) );
  DLH_X1 EK0_temp_expanded_key_reg_127_ ( .G(EK0_n565), .D(EK0_n58), .Q(
        n[3124]) );
  DLH_X1 EK0_temp_expanded_key_reg_95_ ( .G(EK0_n566), .D(EK0_n90), .Q(n[3092]) );
  DLH_X1 EK0_temp_expanded_key_reg_63_ ( .G(EK0_n565), .D(EK0_n122), .Q(
        n[3060]) );
  DLH_X1 EK0_temp_expanded_key_reg_31_ ( .G(EK0_n566), .D(EK0_n154), .Q(
        n[3028]) );
  DFF_X1 EK0_sub_word_reg_31_ ( .D(EK0_n184), .CK(clk), .Q(EK0_n194) );
  DFF_X1 EK0_ready_reg ( .D(EK0_n314), .CK(clk), .Q(n2996) );
  DFF_X1 EK0_cnt_reg_1_ ( .D(EK0_U4_Z_1), .CK(clk), .Q(EK0_add_99_A_1_), .QN(
        EK0_n196) );
  DFF_X1 EK0_cnt_reg_0_ ( .D(EK0_U4_Z_0), .CK(clk), .Q(EK0_add_99_A_0_), .QN(
        EK0_n200) );
  INV_X1 EK0_SB2_U470 ( .A(EK0_SB2_n462), .ZN(EK0_SB2_n461) );
  NOR2_X1 EK0_SB2_U469 ( .A1(EK0_SB2_n89), .A2(EK0_U9_Z_3), .ZN(EK0_SB2_n172)
         );
  NOR2_X1 EK0_SB2_U468 ( .A1(EK0_SB2_n83), .A2(EK0_U9_Z_3), .ZN(EK0_SB2_n133)
         );
  NOR2_X1 EK0_SB2_U467 ( .A1(EK0_SB2_n59), .A2(EK0_U9_Z_3), .ZN(EK0_SB2_n110)
         );
  NOR2_X1 EK0_SB2_U466 ( .A1(EK0_SB2_n50), .A2(EK0_U9_Z_3), .ZN(EK0_SB2_n297)
         );
  AOI211_X1 EK0_SB2_U465 ( .C1(EK0_SB2_n171), .C2(EK0_SB2_n70), .A(
        EK0_SB2_n185), .B(EK0_SB2_n123), .ZN(EK0_SB2_n406) );
  NOR2_X1 EK0_SB2_U460 ( .A1(EK0_U9_Z_3), .A2(EK0_U9_Z_4), .ZN(EK0_SB2_n259)
         );
  NOR2_X1 EK0_SB2_U449 ( .A1(EK0_SB2_n88), .A2(EK0_U9_Z_3), .ZN(EK0_SB2_n454)
         );
  AOI221_X1 EK0_SB2_U445 ( .B1(EK0_SB2_n121), .B2(EK0_SB2_n185), .C1(
        EK0_SB2_n173), .C2(EK0_SB2_n135), .A(EK0_SB2_n46), .ZN(EK0_SB2_n341)
         );
  NOR2_X1 EK0_SB2_U438 ( .A1(EK0_SB2_n18), .A2(EK0_U9_Z_3), .ZN(EK0_SB2_n132)
         );
  AOI22_X1 EK0_SB2_U419 ( .A1(EK0_SB2_n287), .A2(EK0_SB2_n288), .B1(
        EK0_SB2_n89), .B2(EK0_SB2_n185), .ZN(EK0_SB2_n285) );
  AOI21_X1 EK0_SB2_U418 ( .B1(EK0_SB2_n185), .B2(EK0_SB2_n206), .A(
        EK0_SB2_n162), .ZN(EK0_SB2_n182) );
  AOI22_X1 EK0_SB2_U417 ( .A1(EK0_SB2_n190), .A2(EK0_SB2_n298), .B1(
        EK0_SB2_n149), .B2(EK0_SB2_n185), .ZN(EK0_SB2_n353) );
  NOR2_X1 EK0_SB2_U416 ( .A1(EK0_SB2_n185), .A2(EK0_SB2_n157), .ZN(
        EK0_SB2_n230) );
  OAI221_X1 EK0_SB2_U415 ( .B1(EK0_U9_Z_3), .B2(EK0_SB2_n334), .C1(
        EK0_SB2_n439), .C2(EK0_SB2_n35), .A(EK0_SB2_n440), .ZN(EK0_SB2_n433)
         );
  NOR3_X1 EK0_SB2_U414 ( .A1(EK0_SB2_n80), .A2(EK0_U9_Z_3), .A3(EK0_SB2_n28), 
        .ZN(EK0_SB2_n276) );
  OAI22_X1 EK0_SB2_U413 ( .A1(EK0_U9_Z_3), .A2(EK0_SB2_n337), .B1(EK0_SB2_n338), .B2(EK0_SB2_n82), .ZN(EK0_SB2_n336) );
  OAI221_X1 EK0_SB2_U412 ( .B1(EK0_U9_Z_3), .B2(EK0_SB2_n267), .C1(EK0_SB2_n68), .C2(EK0_SB2_n45), .A(EK0_SB2_n268), .ZN(EK0_SB2_n263) );
  AOI222_X1 EK0_SB2_U411 ( .A1(EK0_SB2_n134), .A2(EK0_SB2_n263), .B1(
        EK0_SB2_n264), .B2(EK0_SB2_n185), .C1(EK0_SB2_n133), .C2(EK0_SB2_n265), 
        .ZN(EK0_SB2_n222) );
  OAI22_X1 EK0_SB2_U410 ( .A1(EK0_SB2_n185), .A2(EK0_SB2_n7), .B1(EK0_SB2_n11), 
        .B2(EK0_SB2_n62), .ZN(EK0_SB2_n455) );
  NOR4_X1 EK0_SB2_U409 ( .A1(EK0_SB2_n358), .A2(EK0_SB2_n359), .A3(
        EK0_SB2_n360), .A4(EK0_SB2_n241), .ZN(EK0_SB2_n357) );
  NAND2_X1 EK0_SB2_U408 ( .A1(EK0_SB2_n408), .A2(EK0_SB2_n246), .ZN(
        EK0_SB2_n327) );
  AOI22_X1 EK0_SB2_U407 ( .A1(EK0_SB2_n36), .A2(EK0_SB2_n461), .B1(
        EK0_SB2_n134), .B2(EK0_SB2_n246), .ZN(EK0_SB2_n415) );
  NOR3_X1 EK0_SB2_U406 ( .A1(EK0_SB2_n36), .A2(EK0_SB2_n277), .A3(EK0_SB2_n236), .ZN(EK0_SB2_n449) );
  NAND2_X1 EK0_SB2_U405 ( .A1(EK0_SB2_n137), .A2(EK0_SB2_n246), .ZN(
        EK0_SB2_n342) );
  OAI21_X1 EK0_SB2_U404 ( .B1(EK0_SB2_n235), .B2(EK0_SB2_n236), .A(
        EK0_SB2_n219), .ZN(EK0_SB2_n233) );
  AOI222_X1 EK0_SB2_U403 ( .A1(EK0_SB2_n324), .A2(EK0_SB2_n167), .B1(
        EK0_SB2_n413), .B2(EK0_SB2_n236), .C1(EK0_SB2_n157), .C2(EK0_SB2_n414), 
        .ZN(EK0_SB2_n389) );
  NOR4_X1 EK0_SB2_U402 ( .A1(EK0_SB2_n451), .A2(EK0_SB2_n27), .A3(EK0_SB2_n360), .A4(EK0_SB2_n276), .ZN(EK0_SB2_n429) );
  OAI221_X1 EK0_SB2_U401 ( .B1(EK0_SB2_n321), .B2(EK0_SB2_n54), .C1(
        EK0_SB2_n322), .C2(EK0_SB2_n64), .A(EK0_SB2_n323), .ZN(EK0_SB2_n319)
         );
  INV_X1 EK0_SB2_U400 ( .A(EK0_n569), .ZN(EK0_SB2_n41) );
  AOI221_X1 EK0_SB2_U399 ( .B1(EK0_SB2_n123), .B2(EK0_SB2_n370), .C1(
        EK0_SB2_n162), .C2(EK0_SB2_n124), .A(EK0_SB2_n371), .ZN(EK0_SB2_n355)
         );
  OAI222_X1 EK0_SB2_U398 ( .A1(EK0_SB2_n284), .A2(EK0_SB2_n56), .B1(
        EK0_SB2_n285), .B2(EK0_SB2_n38), .C1(EK0_SB2_n459), .C2(EK0_SB2_n286), 
        .ZN(EK0_SB2_n283) );
  NOR3_X1 EK0_SB2_U397 ( .A1(EK0_SB2_n301), .A2(EK0_SB2_n193), .A3(
        EK0_SB2_n302), .ZN(EK0_SB2_n292) );
  OAI222_X1 EK0_SB2_U396 ( .A1(EK0_SB2_n292), .A2(EK0_SB2_n62), .B1(
        EK0_SB2_n293), .B2(EK0_SB2_n30), .C1(EK0_SB2_n294), .C2(EK0_SB2_n7), 
        .ZN(EK0_SB2_n291) );
  INV_X1 EK0_SB2_U395 ( .A(EK0_U9_Z_1), .ZN(EK0_SB2_n460) );
  INV_X1 EK0_SB2_U394 ( .A(EK0_U9_Z_0), .ZN(EK0_SB2_n462) );
  AOI22_X1 EK0_SB2_U393 ( .A1(EK0_SB2_n136), .A2(EK0_SB2_n155), .B1(
        EK0_SB2_n36), .B2(EK0_SB2_n123), .ZN(EK0_SB2_n154) );
  OAI21_X1 EK0_SB2_U392 ( .B1(EK0_SB2_n156), .B2(EK0_SB2_n12), .A(EK0_SB2_n157), .ZN(EK0_SB2_n152) );
  NOR2_X1 EK0_SB2_U391 ( .A1(EK0_n286), .A2(EK0_SB2_n50), .ZN(EK0_SB2_n380) );
  OAI22_X1 EK0_SB2_U390 ( .A1(EK0_n286), .A2(EK0_SB2_n37), .B1(EK0_SB2_n55), 
        .B2(EK0_SB2_n11), .ZN(EK0_SB2_n155) );
  OAI22_X1 EK0_SB2_U389 ( .A1(EK0_SB2_n84), .A2(EK0_SB2_n66), .B1(EK0_SB2_n68), 
        .B2(EK0_SB2_n88), .ZN(EK0_SB2_n201) );
  NOR2_X1 EK0_SB2_U388 ( .A1(EK0_SB2_n45), .A2(EK0_n286), .ZN(EK0_SB2_n235) );
  NOR3_X1 EK0_SB2_U387 ( .A1(EK0_SB2_n50), .A2(EK0_n286), .A3(EK0_SB2_n101), 
        .ZN(EK0_SB2_n118) );
  OAI21_X1 EK0_SB2_U386 ( .B1(EK0_SB2_n37), .B2(EK0_SB2_n60), .A(EK0_SB2_n4), 
        .ZN(EK0_SB2_n252) );
  OAI211_X1 EK0_SB2_U385 ( .C1(EK0_SB2_n452), .C2(EK0_SB2_n65), .A(EK0_SB2_n53), .B(EK0_SB2_n60), .ZN(EK0_SB2_n253) );
  AOI221_X1 EK0_SB2_U384 ( .B1(EK0_SB2_n136), .B2(EK0_SB2_n252), .C1(
        EK0_SB2_n213), .C2(EK0_SB2_n253), .A(EK0_SB2_n254), .ZN(EK0_SB2_n251)
         );
  OAI21_X1 EK0_SB2_U383 ( .B1(EK0_SB2_n49), .B2(EK0_SB2_n35), .A(EK0_SB2_n19), 
        .ZN(EK0_SB2_n425) );
  NOR2_X1 EK0_SB2_U382 ( .A1(EK0_n286), .A2(EK0_U9_Z_4), .ZN(EK0_SB2_n426) );
  AOI221_X1 EK0_SB2_U381 ( .B1(EK0_SB2_n136), .B2(EK0_SB2_n425), .C1(
        EK0_SB2_n426), .C2(EK0_SB2_n133), .A(EK0_SB2_n159), .ZN(EK0_SB2_n424)
         );
  NOR2_X1 EK0_SB2_U380 ( .A1(EK0_SB2_n452), .A2(EK0_n286), .ZN(EK0_SB2_n206)
         );
  NOR3_X1 EK0_SB2_U379 ( .A1(EK0_SB2_n64), .A2(EK0_n286), .A3(EK0_SB2_n59), 
        .ZN(EK0_SB2_n310) );
  OAI22_X1 EK0_SB2_U378 ( .A1(EK0_n569), .A2(EK0_U9_Z_4), .B1(EK0_SB2_n452), 
        .B2(EK0_SB2_n30), .ZN(EK0_SB2_n309) );
  AOI221_X1 EK0_SB2_U377 ( .B1(EK0_SB2_n160), .B2(EK0_SB2_n124), .C1(
        EK0_SB2_n157), .C2(EK0_SB2_n309), .A(EK0_SB2_n310), .ZN(EK0_SB2_n308)
         );
  NOR2_X1 EK0_SB2_U376 ( .A1(EK0_n569), .A2(EK0_n286), .ZN(EK0_SB2_n213) );
  NAND2_X1 EK0_SB2_U375 ( .A1(EK0_SB2_n172), .A2(EK0_n286), .ZN(EK0_SB2_n443)
         );
  NAND2_X1 EK0_SB2_U374 ( .A1(EK0_SB2_n459), .A2(EK0_n569), .ZN(EK0_SB2_n210)
         );
  NAND2_X1 EK0_SB2_U373 ( .A1(EK0_SB2_n235), .A2(EK0_SB2_n105), .ZN(
        EK0_SB2_n334) );
  NAND2_X1 EK0_SB2_U372 ( .A1(EK0_SB2_n245), .A2(EK0_SB2_n32), .ZN(
        EK0_SB2_n142) );
  NAND2_X1 EK0_SB2_U371 ( .A1(EK0_SB2_n452), .A2(EK0_SB2_n41), .ZN(
        EK0_SB2_n145) );
  OAI21_X1 EK0_SB2_U370 ( .B1(EK0_SB2_n140), .B2(EK0_SB2_n141), .A(
        EK0_SB2_n142), .ZN(EK0_SB2_n139) );
  INV_X1 EK0_SB2_U369 ( .A(EK0_SB2_n139), .ZN(EK0_SB2_n26) );
  OAI211_X1 EK0_SB2_U368 ( .C1(EK0_SB2_n18), .C2(EK0_SB2_n65), .A(EK0_SB2_n138), .B(EK0_SB2_n26), .ZN(EK0_SB2_n128) );
  NAND2_X1 EK0_SB2_U367 ( .A1(EK0_SB2_n89), .A2(EK0_SB2_n452), .ZN(
        EK0_SB2_n307) );
  AOI21_X1 EK0_SB2_U366 ( .B1(EK0_SB2_n64), .B2(EK0_SB2_n307), .A(EK0_SB2_n35), 
        .ZN(EK0_SB2_n387) );
  AOI211_X1 EK0_SB2_U365 ( .C1(EK0_SB2_n386), .C2(EK0_SB2_n83), .A(
        EK0_SB2_n282), .B(EK0_SB2_n387), .ZN(EK0_SB2_n385) );
  AOI22_X1 EK0_SB2_U364 ( .A1(EK0_SB2_n235), .A2(EK0_SB2_n70), .B1(
        EK0_SB2_n237), .B2(EK0_SB2_n143), .ZN(EK0_SB2_n384) );
  OAI211_X1 EK0_SB2_U363 ( .C1(EK0_SB2_n7), .C2(EK0_SB2_n49), .A(EK0_SB2_n384), 
        .B(EK0_SB2_n385), .ZN(EK0_SB2_n382) );
  OAI21_X1 EK0_SB2_U362 ( .B1(EK0_SB2_n58), .B2(EK0_SB2_n84), .A(EK0_SB2_n170), 
        .ZN(EK0_SB2_n169) );
  AOI221_X1 EK0_SB2_U361 ( .B1(EK0_SB2_n110), .B2(EK0_SB2_n167), .C1(
        EK0_SB2_n168), .C2(EK0_SB2_n135), .A(EK0_SB2_n169), .ZN(EK0_SB2_n166)
         );
  AOI22_X1 EK0_SB2_U360 ( .A1(EK0_SB2_n173), .A2(EK0_SB2_n452), .B1(
        EK0_SB2_n137), .B2(EK0_SB2_n144), .ZN(EK0_SB2_n165) );
  OAI211_X1 EK0_SB2_U359 ( .C1(EK0_SB2_n85), .C2(EK0_SB2_n66), .A(EK0_SB2_n165), .B(EK0_SB2_n166), .ZN(EK0_SB2_n164) );
  NOR3_X1 EK0_SB2_U358 ( .A1(EK0_SB2_n63), .A2(EK0_U9_Z_4), .A3(EK0_SB2_n32), 
        .ZN(EK0_SB2_n359) );
  NOR2_X1 EK0_SB2_U357 ( .A1(EK0_SB2_n452), .A2(EK0_SB2_n83), .ZN(EK0_SB2_n191) );
  AOI22_X1 EK0_SB2_U356 ( .A1(EK0_SB2_n191), .A2(EK0_SB2_n105), .B1(
        EK0_SB2_n171), .B2(EK0_SB2_n192), .ZN(EK0_SB2_n189) );
  AOI221_X1 EK0_SB2_U355 ( .B1(EK0_SB2_n105), .B2(EK0_SB2_n382), .C1(
        EK0_SB2_n350), .C2(EK0_SB2_n453), .A(EK0_SB2_n383), .ZN(EK0_SB2_n354)
         );
  AOI221_X1 EK0_SB2_U354 ( .B1(EK0_SB2_n163), .B2(EK0_SB2_n361), .C1(
        EK0_SB2_n213), .C2(EK0_SB2_n362), .A(EK0_SB2_n363), .ZN(EK0_SB2_n356)
         );
  NAND4_X1 EK0_SB2_U353 ( .A1(EK0_SB2_n354), .A2(EK0_SB2_n355), .A3(
        EK0_SB2_n356), .A4(EK0_SB2_n357), .ZN(EK0_n280) );
  AOI221_X1 EK0_SB2_U352 ( .B1(EK0_SB2_n350), .B2(EK0_SB2_n149), .C1(
        EK0_SB2_n156), .C2(EK0_SB2_n124), .A(EK0_SB2_n402), .ZN(EK0_SB2_n390)
         );
  NOR4_X1 EK0_SB2_U351 ( .A1(EK0_SB2_n392), .A2(EK0_SB2_n393), .A3(
        EK0_SB2_n394), .A4(EK0_SB2_n395), .ZN(EK0_SB2_n391) );
  NAND4_X1 EK0_SB2_U350 ( .A1(EK0_SB2_n388), .A2(EK0_SB2_n389), .A3(
        EK0_SB2_n390), .A4(EK0_SB2_n391), .ZN(EK0_n279) );
  NAND2_X1 EK0_SB2_U349 ( .A1(EK0_SB2_n163), .A2(EK0_SB2_n408), .ZN(
        EK0_SB2_n113) );
  AOI22_X1 EK0_SB2_U348 ( .A1(EK0_SB2_n237), .A2(EK0_SB2_n148), .B1(
        EK0_SB2_n12), .B2(EK0_SB2_n70), .ZN(EK0_SB2_n232) );
  OAI21_X1 EK0_SB2_U347 ( .B1(EK0_SB2_n121), .B2(EK0_SB2_n124), .A(EK0_SB2_n31), .ZN(EK0_SB2_n234) );
  OAI211_X1 EK0_SB2_U346 ( .C1(EK0_SB2_n232), .C2(EK0_SB2_n84), .A(
        EK0_SB2_n233), .B(EK0_SB2_n234), .ZN(EK0_SB2_n227) );
  AOI221_X1 EK0_SB2_U345 ( .B1(EK0_SB2_n31), .B2(EK0_SB2_n123), .C1(
        EK0_SB2_n288), .C2(EK0_SB2_n213), .A(EK0_SB2_n217), .ZN(EK0_SB2_n332)
         );
  INV_X1 EK0_SB2_U344 ( .A(EK0_SB2_n282), .ZN(EK0_SB2_n22) );
  OAI22_X1 EK0_SB2_U343 ( .A1(EK0_SB2_n332), .A2(EK0_SB2_n88), .B1(EK0_SB2_n75), .B2(EK0_SB2_n22), .ZN(EK0_SB2_n331) );
  INV_X1 EK0_SB2_U342 ( .A(EK0_SB2_n89), .ZN(EK0_SB2_n83) );
  OAI22_X1 EK0_SB2_U341 ( .A1(EK0_SB2_n460), .A2(EK0_SB2_n15), .B1(
        EK0_SB2_n287), .B2(EK0_SB2_n5), .ZN(EK0_SB2_n301) );
  NOR3_X1 EK0_SB2_U340 ( .A1(EK0_SB2_n23), .A2(EK0_SB2_n452), .A3(EK0_SB2_n453), .ZN(EK0_SB2_n302) );
  NOR4_X1 EK0_SB2_U339 ( .A1(EK0_SB2_n226), .A2(EK0_SB2_n227), .A3(
        EK0_SB2_n228), .A4(EK0_SB2_n229), .ZN(EK0_SB2_n225) );
  AOI221_X1 EK0_SB2_U338 ( .B1(EK0_SB2_n120), .B2(EK0_SB2_n260), .C1(
        EK0_SB2_n213), .C2(EK0_SB2_n261), .A(EK0_SB2_n262), .ZN(EK0_SB2_n223)
         );
  NOR2_X1 EK0_SB2_U337 ( .A1(EK0_U9_Z_4), .A2(EK0_SB2_n452), .ZN(EK0_SB2_n298)
         );
  INV_X1 EK0_SB2_U336 ( .A(EK0_SB2_n452), .ZN(EK0_SB2_n50) );
  OAI222_X1 EK0_SB2_U335 ( .A1(EK0_SB2_n197), .A2(EK0_SB2_n5), .B1(EK0_U9_Z_0), 
        .B2(EK0_SB2_n251), .C1(EK0_SB2_n81), .C2(EK0_SB2_n113), .ZN(
        EK0_SB2_n248) );
  OAI22_X1 EK0_SB2_U334 ( .A1(EK0_SB2_n250), .A2(EK0_SB2_n21), .B1(EK0_SB2_n72), .B2(EK0_SB2_n114), .ZN(EK0_SB2_n249) );
  AOI211_X1 EK0_SB2_U333 ( .C1(EK0_SB2_n163), .C2(EK0_SB2_n247), .A(
        EK0_SB2_n248), .B(EK0_SB2_n249), .ZN(EK0_SB2_n224) );
  OAI211_X1 EK0_SB2_U332 ( .C1(EK0_SB2_n194), .C2(EK0_SB2_n88), .A(
        EK0_SB2_n195), .B(EK0_SB2_n196), .ZN(EK0_SB2_n179) );
  OAI222_X1 EK0_SB2_U331 ( .A1(EK0_SB2_n64), .A2(EK0_SB2_n17), .B1(
        EK0_SB2_n189), .B2(EK0_SB2_n35), .C1(EK0_SB2_n67), .C2(EK0_SB2_n2), 
        .ZN(EK0_SB2_n180) );
  NOR4_X1 EK0_SB2_U330 ( .A1(EK0_SB2_n178), .A2(EK0_SB2_n179), .A3(
        EK0_SB2_n180), .A4(EK0_SB2_n181), .ZN(EK0_SB2_n177) );
  NOR2_X1 EK0_SB2_U329 ( .A1(EK0_SB2_n89), .A2(EK0_U9_Z_4), .ZN(EK0_SB2_n269)
         );
  AOI222_X1 EK0_SB2_U328 ( .A1(EK0_SB2_n126), .A2(EK0_SB2_n143), .B1(
        EK0_SB2_n269), .B2(EK0_SB2_n102), .C1(EK0_SB2_n206), .C2(EK0_SB2_n104), 
        .ZN(EK0_SB2_n268) );
  AOI22_X1 EK0_SB2_U327 ( .A1(EK0_SB2_n89), .A2(EK0_SB2_n277), .B1(
        EK0_SB2_n120), .B2(EK0_SB2_n202), .ZN(EK0_SB2_n204) );
  NOR2_X1 EK0_SB2_U326 ( .A1(EK0_SB2_n59), .A2(EK0_SB2_n89), .ZN(EK0_SB2_n104)
         );
  AOI21_X1 EK0_SB2_U325 ( .B1(EK0_SB2_n134), .B2(EK0_SB2_n368), .A(EK0_SB2_n1), 
        .ZN(EK0_SB2_n364) );
  AND3_X1 EK0_SB2_U324 ( .A1(EK0_SB2_n367), .A2(EK0_SB2_n75), .A3(EK0_SB2_n64), 
        .ZN(EK0_SB2_n365) );
  INV_X1 EK0_SB2_U323 ( .A(EK0_SB2_n366), .ZN(EK0_SB2_n10) );
  OAI221_X1 EK0_SB2_U322 ( .B1(EK0_SB2_n89), .B2(EK0_SB2_n364), .C1(
        EK0_SB2_n365), .C2(EK0_SB2_n2), .A(EK0_SB2_n10), .ZN(EK0_SB2_n363) );
  NOR2_X1 EK0_SB2_U321 ( .A1(EK0_SB2_n59), .A2(EK0_SB2_n452), .ZN(EK0_SB2_n221) );
  AOI22_X1 EK0_SB2_U320 ( .A1(EK0_SB2_n117), .A2(EK0_SB2_n288), .B1(
        EK0_SB2_n172), .B2(EK0_SB2_n163), .ZN(EK0_SB2_n348) );
  AOI21_X1 EK0_SB2_U319 ( .B1(EK0_SB2_n59), .B2(EK0_SB2_n32), .A(EK0_SB2_n148), 
        .ZN(EK0_SB2_n438) );
  OAI222_X1 EK0_SB2_U318 ( .A1(EK0_SB2_n70), .A2(EK0_SB2_n28), .B1(
        EK0_SB2_n438), .B2(EK0_SB2_n68), .C1(EK0_SB2_n49), .C2(EK0_SB2_n35), 
        .ZN(EK0_SB2_n436) );
  OAI22_X1 EK0_SB2_U317 ( .A1(EK0_SB2_n64), .A2(EK0_SB2_n267), .B1(EK0_SB2_n51), .B2(EK0_SB2_n69), .ZN(EK0_SB2_n437) );
  AOI211_X1 EK0_SB2_U316 ( .C1(EK0_SB2_n124), .C2(EK0_SB2_n103), .A(
        EK0_SB2_n436), .B(EK0_SB2_n437), .ZN(EK0_SB2_n435) );
  NOR3_X1 EK0_SB2_U315 ( .A1(EK0_SB2_n73), .A2(EK0_n569), .A3(EK0_SB2_n44), 
        .ZN(EK0_SB2_n340) );
  AOI211_X1 EK0_SB2_U314 ( .C1(EK0_SB2_n126), .C2(EK0_SB2_n103), .A(
        EK0_SB2_n31), .B(EK0_SB2_n188), .ZN(EK0_SB2_n338) );
  AOI221_X1 EK0_SB2_U312 ( .B1(EK0_SB2_n324), .B2(EK0_SB2_n462), .C1(
        EK0_SB2_n339), .C2(EK0_SB2_n231), .A(EK0_SB2_n340), .ZN(EK0_SB2_n337)
         );
  AOI221_X1 EK0_SB2_U311 ( .B1(EK0_SB2_n126), .B2(EK0_SB2_n127), .C1(
        EK0_SB2_n461), .C2(EK0_SB2_n128), .A(EK0_SB2_n129), .ZN(EK0_SB2_n92)
         );
  AOI22_X1 EK0_SB2_U310 ( .A1(EK0_SB2_n162), .A2(EK0_SB2_n144), .B1(
        EK0_SB2_n163), .B2(EK0_SB2_n164), .ZN(EK0_SB2_n90) );
  AOI22_X1 EK0_SB2_U309 ( .A1(EK0_SB2_n459), .A2(EK0_SB2_n150), .B1(
        EK0_SB2_n151), .B2(EK0_SB2_n462), .ZN(EK0_SB2_n91) );
  AOI221_X1 EK0_SB2_U308 ( .B1(EK0_SB2_n143), .B2(EK0_SB2_n343), .C1(
        EK0_SB2_n162), .C2(EK0_SB2_n157), .A(EK0_SB2_n344), .ZN(EK0_SB2_n314)
         );
  AOI221_X1 EK0_SB2_U307 ( .B1(EK0_SB2_n24), .B2(EK0_SB2_n219), .C1(
        EK0_SB2_n163), .C2(EK0_SB2_n335), .A(EK0_SB2_n336), .ZN(EK0_SB2_n315)
         );
  AOI221_X1 EK0_SB2_U306 ( .B1(EK0_SB2_n89), .B2(EK0_SB2_n329), .C1(
        EK0_SB2_n160), .C2(EK0_SB2_n330), .A(EK0_SB2_n331), .ZN(EK0_SB2_n316)
         );
  AOI211_X1 EK0_SB2_U305 ( .C1(EK0_SB2_n202), .C2(EK0_SB2_n157), .A(
        EK0_SB2_n203), .B(EK0_SB2_n3), .ZN(EK0_SB2_n176) );
  AOI222_X1 EK0_SB2_U304 ( .A1(EK0_SB2_n143), .A2(EK0_SB2_n211), .B1(
        EK0_SB2_n31), .B2(EK0_SB2_n212), .C1(EK0_SB2_n213), .C2(EK0_SB2_n214), 
        .ZN(EK0_SB2_n175) );
  AOI222_X1 EK0_SB2_U303 ( .A1(EK0_SB2_n144), .A2(EK0_SB2_n217), .B1(
        EK0_SB2_n134), .B2(EK0_SB2_n218), .C1(EK0_SB2_n219), .C2(EK0_SB2_n40), 
        .ZN(EK0_SB2_n174) );
  AOI221_X1 EK0_SB2_U302 ( .B1(EK0_SB2_n109), .B2(EK0_SB2_n460), .C1(
        EK0_SB2_n110), .C2(EK0_SB2_n111), .A(EK0_SB2_n112), .ZN(EK0_SB2_n108)
         );
  AOI211_X1 EK0_SB2_U301 ( .C1(EK0_SB2_n116), .C2(EK0_SB2_n117), .A(
        EK0_SB2_n118), .B(EK0_SB2_n119), .ZN(EK0_SB2_n107) );
  AOI22_X1 EK0_SB2_U300 ( .A1(EK0_SB2_n122), .A2(EK0_SB2_n123), .B1(
        EK0_SB2_n124), .B2(EK0_SB2_n125), .ZN(EK0_SB2_n106) );
  OAI221_X1 EK0_SB2_U299 ( .B1(EK0_n569), .B2(EK0_SB2_n106), .C1(EK0_SB2_n107), 
        .C2(EK0_SB2_n54), .A(EK0_SB2_n108), .ZN(EK0_SB2_n94) );
  NOR2_X1 EK0_SB2_U298 ( .A1(EK0_SB2_n83), .A2(EK0_U9_Z_4), .ZN(EK0_SB2_n237)
         );
  NOR2_X1 EK0_SB2_U297 ( .A1(EK0_SB2_n32), .A2(EK0_SB2_n50), .ZN(EK0_SB2_n281)
         );
  OAI221_X1 EK0_SB2_U296 ( .B1(EK0_SB2_n9), .B2(EK0_SB2_n69), .C1(EK0_SB2_n65), 
        .C2(EK0_SB2_n2), .A(EK0_SB2_n308), .ZN(EK0_SB2_n289) );
  OAI211_X1 EK0_SB2_U295 ( .C1(EK0_SB2_n56), .C2(EK0_SB2_n82), .A(EK0_SB2_n303), .B(EK0_SB2_n304), .ZN(EK0_SB2_n290) );
  AOI221_X1 EK0_SB2_U294 ( .B1(EK0_U9_Z_0), .B2(EK0_SB2_n289), .C1(
        EK0_SB2_n163), .C2(EK0_SB2_n290), .A(EK0_SB2_n291), .ZN(EK0_SB2_n271)
         );
  AOI21_X1 EK0_SB2_U293 ( .B1(EK0_SB2_n78), .B2(EK0_SB2_n76), .A(EK0_SB2_n54), 
        .ZN(EK0_SB2_n441) );
  AOI221_X1 EK0_SB2_U292 ( .B1(EK0_SB2_n171), .B2(EK0_SB2_n444), .C1(
        EK0_SB2_n445), .C2(EK0_SB2_n50), .A(EK0_SB2_n446), .ZN(EK0_SB2_n439)
         );
  OAI21_X1 EK0_SB2_U291 ( .B1(EK0_SB2_n441), .B2(EK0_SB2_n442), .A(
        EK0_SB2_n102), .ZN(EK0_SB2_n440) );
  AOI222_X1 EK0_SB2_U290 ( .A1(EK0_SB2_n173), .A2(EK0_SB2_n452), .B1(
        EK0_SB2_n137), .B2(EK0_SB2_n167), .C1(EK0_SB2_n168), .C2(EK0_SB2_n259), 
        .ZN(EK0_SB2_n258) );
  NOR2_X1 EK0_SB2_U289 ( .A1(EK0_SB2_n461), .A2(EK0_SB2_n89), .ZN(EK0_SB2_n121) );
  OAI222_X1 EK0_SB2_U288 ( .A1(EK0_SB2_n459), .A2(EK0_SB2_n38), .B1(
        EK0_SB2_n30), .B2(EK0_SB2_n88), .C1(EK0_SB2_n7), .C2(EK0_SB2_n82), 
        .ZN(EK0_SB2_n208) );
  AOI211_X1 EK0_SB2_U287 ( .C1(EK0_SB2_n206), .C2(EK0_SB2_n207), .A(
        EK0_SB2_n208), .B(EK0_SB2_n209), .ZN(EK0_SB2_n205) );
  OAI222_X1 EK0_SB2_U286 ( .A1(EK0_SB2_n80), .A2(EK0_SB2_n15), .B1(
        EK0_SB2_n205), .B2(EK0_SB2_n54), .C1(EK0_SB2_n81), .C2(EK0_SB2_n115), 
        .ZN(EK0_SB2_n203) );
  OAI211_X1 EK0_SB2_U285 ( .C1(EK0_SB2_n34), .C2(EK0_SB2_n69), .A(EK0_SB2_n204), .B(EK0_SB2_n424), .ZN(EK0_SB2_n416) );
  OAI221_X1 EK0_SB2_U284 ( .B1(EK0_SB2_n43), .B2(EK0_SB2_n75), .C1(EK0_SB2_n73), .C2(EK0_SB2_n45), .A(EK0_SB2_n419), .ZN(EK0_SB2_n418) );
  AOI222_X1 EK0_SB2_U283 ( .A1(EK0_SB2_n416), .A2(EK0_SB2_n462), .B1(
        EK0_SB2_n417), .B2(EK0_SB2_n59), .C1(EK0_SB2_n163), .C2(EK0_SB2_n418), 
        .ZN(EK0_SB2_n388) );
  NOR3_X1 EK0_SB2_U282 ( .A1(EK0_SB2_n11), .A2(EK0_n569), .A3(EK0_SB2_n70), 
        .ZN(EK0_SB2_n186) );
  AOI211_X1 EK0_SB2_U281 ( .C1(EK0_SB2_n163), .C2(EK0_SB2_n185), .A(
        EK0_SB2_n156), .B(EK0_SB2_n186), .ZN(EK0_SB2_n184) );
  AOI221_X1 EK0_SB2_U280 ( .B1(EK0_SB2_n110), .B2(EK0_SB2_n102), .C1(
        EK0_SB2_n126), .C2(EK0_SB2_n187), .A(EK0_SB2_n188), .ZN(EK0_SB2_n183)
         );
  OAI222_X1 EK0_SB2_U279 ( .A1(EK0_SB2_n182), .A2(EK0_SB2_n74), .B1(
        EK0_SB2_n183), .B2(EK0_SB2_n76), .C1(EK0_SB2_n184), .C2(EK0_SB2_n78), 
        .ZN(EK0_SB2_n181) );
  AOI21_X1 EK0_SB2_U278 ( .B1(EK0_SB2_n160), .B2(EK0_SB2_n157), .A(
        EK0_SB2_n159), .ZN(EK0_SB2_n286) );
  AOI22_X1 EK0_SB2_U277 ( .A1(EK0_SB2_n117), .A2(EK0_SB2_n207), .B1(
        EK0_SB2_n120), .B2(EK0_SB2_n148), .ZN(EK0_SB2_n284) );
  INV_X1 EK0_SB2_U276 ( .A(EK0_SB2_n213), .ZN(EK0_SB2_n7) );
  NOR2_X1 EK0_SB2_U275 ( .A1(EK0_SB2_n41), .A2(EK0_SB2_n452), .ZN(EK0_SB2_n148) );
  AOI221_X1 EK0_SB2_U274 ( .B1(EK0_SB2_n231), .B2(EK0_SB2_n379), .C1(
        EK0_SB2_n380), .C2(EK0_SB2_n287), .A(EK0_SB2_n381), .ZN(EK0_SB2_n378)
         );
  OAI222_X1 EK0_SB2_U273 ( .A1(EK0_SB2_n372), .A2(EK0_SB2_n66), .B1(
        EK0_SB2_n78), .B2(EK0_SB2_n342), .C1(EK0_SB2_n373), .C2(EK0_SB2_n30), 
        .ZN(EK0_SB2_n371) );
  OAI221_X1 EK0_SB2_U272 ( .B1(EK0_SB2_n460), .B2(EK0_SB2_n327), .C1(
        EK0_SB2_n461), .C2(EK0_SB2_n2), .A(EK0_SB2_n378), .ZN(EK0_SB2_n370) );
  NOR2_X1 EK0_SB2_U271 ( .A1(EK0_SB2_n70), .A2(EK0_SB2_n89), .ZN(EK0_SB2_n123)
         );
  NOR2_X1 EK0_SB2_U270 ( .A1(EK0_SB2_n452), .A2(EK0_n569), .ZN(EK0_SB2_n102)
         );
  NOR2_X1 EK0_SB2_U269 ( .A1(EK0_SB2_n462), .A2(EK0_SB2_n89), .ZN(EK0_SB2_n219) );
  NOR2_X1 EK0_SB2_U268 ( .A1(EK0_SB2_n32), .A2(EK0_SB2_n452), .ZN(EK0_SB2_n117) );
  NOR2_X1 EK0_SB2_U267 ( .A1(EK0_SB2_n460), .A2(EK0_SB2_n89), .ZN(EK0_SB2_n124) );
  INV_X1 EK0_SB2_U266 ( .A(EK0_SB2_n104), .ZN(EK0_SB2_n58) );
  INV_X1 EK0_SB2_U265 ( .A(EK0_SB2_n204), .ZN(EK0_SB2_n3) );
  OAI222_X1 EK0_SB2_U262 ( .A1(EK0_SB2_n60), .A2(EK0_SB2_n84), .B1(
        EK0_SB2_n307), .B2(EK0_SB2_n88), .C1(EK0_SB2_n43), .C2(EK0_SB2_n82), 
        .ZN(EK0_SB2_n450) );
  INV_X1 EK0_SB2_U261 ( .A(EK0_SB2_n450), .ZN(EK0_SB2_n42) );
  INV_X1 EK0_SB2_U260 ( .A(EK0_SB2_n333), .ZN(EK0_SB2_n1) );
  OR3_X1 EK0_SB2_U259 ( .A1(EK0_SB2_n197), .A2(EK0_SB2_n461), .A3(EK0_SB2_n113), .ZN(EK0_SB2_n195) );
  INV_X1 EK0_SB2_U258 ( .A(EK0_SB2_n237), .ZN(EK0_SB2_n53) );
  AND3_X1 EK0_SB2_U257 ( .A1(EK0_SB2_n136), .A2(EK0_SB2_n103), .A3(
        EK0_SB2_n259), .ZN(EK0_SB2_n87) );
  NOR3_X1 EK0_SB2_U256 ( .A1(EK0_SB2_n55), .A2(EK0_SB2_n250), .A3(EK0_SB2_n23), 
        .ZN(EK0_SB2_n13) );
  OR3_X1 EK0_SB2_U255 ( .A1(EK0_SB2_n13), .A2(EK0_SB2_n240), .A3(EK0_SB2_n87), 
        .ZN(EK0_SB2_n451) );
  INV_X1 EK0_SB2_U254 ( .A(EK0_SB2_n454), .ZN(EK0_SB2_n71) );
  NAND2_X1 EK0_SB2_U253 ( .A1(EK0_SB2_n237), .A2(EK0_SB2_n134), .ZN(
        EK0_SB2_n300) );
  NAND2_X1 EK0_SB2_U252 ( .A1(EK0_SB2_n461), .A2(EK0_SB2_n70), .ZN(
        EK0_SB2_n367) );
  NAND2_X1 EK0_SB2_U251 ( .A1(EK0_SB2_n245), .A2(EK0_SB2_n41), .ZN(
        EK0_SB2_n114) );
  OAI211_X1 EK0_SB2_U250 ( .C1(EK0_SB2_n460), .C2(EK0_SB2_n20), .A(EK0_SB2_n5), 
        .B(EK0_SB2_n415), .ZN(EK0_SB2_n414) );
  OAI211_X1 EK0_SB2_U249 ( .C1(EK0_SB2_n102), .C2(EK0_SB2_n103), .A(
        EK0_SB2_n104), .B(EK0_SB2_n105), .ZN(EK0_SB2_n98) );
  NOR2_X1 EK0_SB2_U248 ( .A1(EK0_SB2_n59), .A2(EK0_SB2_n86), .ZN(EK0_SB2_n122)
         );
  INV_X1 EK0_SB2_U247 ( .A(EK0_SB2_n135), .ZN(EK0_SB2_n43) );
  NAND2_X1 EK0_SB2_U246 ( .A1(EK0_SB2_n124), .A2(EK0_SB2_n143), .ZN(
        EK0_SB2_n140) );
  OAI21_X1 EK0_SB2_U245 ( .B1(EK0_SB2_n7), .B2(EK0_SB2_n54), .A(EK0_SB2_n18), 
        .ZN(EK0_SB2_n386) );
  OAI221_X1 EK0_SB2_U244 ( .B1(EK0_SB2_n64), .B2(EK0_SB2_n145), .C1(
        EK0_SB2_n30), .C2(EK0_SB2_n307), .A(EK0_SB2_n348), .ZN(EK0_SB2_n347)
         );
  OAI21_X1 EK0_SB2_U243 ( .B1(EK0_SB2_n346), .B2(EK0_SB2_n347), .A(
        EK0_SB2_n134), .ZN(EK0_SB2_n345) );
  OAI21_X1 EK0_SB2_U242 ( .B1(EK0_SB2_n74), .B2(EK0_SB2_n21), .A(EK0_SB2_n345), 
        .ZN(EK0_SB2_n344) );
  NAND2_X1 EK0_SB2_U241 ( .A1(EK0_SB2_n287), .A2(EK0_SB2_n281), .ZN(
        EK0_SB2_n146) );
  OAI21_X1 EK0_SB2_U240 ( .B1(EK0_SB2_n168), .B2(EK0_SB2_n70), .A(EK0_SB2_n156), .ZN(EK0_SB2_n196) );
  INV_X1 EK0_SB2_U239 ( .A(EK0_SB2_n219), .ZN(EK0_SB2_n77) );
  INV_X1 EK0_SB2_U238 ( .A(EK0_SB2_n171), .ZN(EK0_SB2_n45) );
  NOR2_X1 EK0_SB2_U237 ( .A1(EK0_SB2_n145), .A2(EK0_SB2_n80), .ZN(EK0_SB2_n264) );
  INV_X1 EK0_SB2_U236 ( .A(EK0_SB2_n281), .ZN(EK0_SB2_n9) );
  NAND2_X1 EK0_SB2_U235 ( .A1(EK0_SB2_n70), .A2(EK0_SB2_n50), .ZN(EK0_SB2_n141) );
  NAND2_X1 EK0_SB2_U234 ( .A1(EK0_SB2_n7), .A2(EK0_SB2_n38), .ZN(EK0_SB2_n326)
         );
  AOI22_X1 EK0_SB2_U233 ( .A1(EK0_SB2_n105), .A2(EK0_SB2_n326), .B1(
        EK0_SB2_n117), .B2(EK0_SB2_n192), .ZN(EK0_SB2_n321) );
  INV_X1 EK0_SB2_U232 ( .A(EK0_SB2_n117), .ZN(EK0_SB2_n11) );
  NOR2_X1 EK0_SB2_U231 ( .A1(EK0_SB2_n64), .A2(EK0_SB2_n460), .ZN(EK0_SB2_n413) );
  AOI21_X1 EK0_SB2_U230 ( .B1(EK0_SB2_n126), .B2(EK0_SB2_n117), .A(
        EK0_SB2_n132), .ZN(EK0_SB2_n194) );
  NAND2_X1 EK0_SB2_U229 ( .A1(EK0_SB2_n143), .A2(EK0_SB2_n231), .ZN(
        EK0_SB2_n130) );
  INV_X1 EK0_SB2_U228 ( .A(EK0_SB2_n460), .ZN(EK0_SB2_n459) );
  AOI21_X1 EK0_SB2_U227 ( .B1(EK0_SB2_n161), .B2(EK0_SB2_n157), .A(
        EK0_SB2_n448), .ZN(EK0_SB2_n447) );
  INV_X1 EK0_SB2_U226 ( .A(EK0_SB2_n113), .ZN(EK0_SB2_n36) );
  NOR2_X1 EK0_SB2_U225 ( .A1(EK0_SB2_n70), .A2(EK0_SB2_n453), .ZN(EK0_SB2_n311) );
  OAI211_X1 EK0_SB2_U224 ( .C1(EK0_SB2_n461), .C2(EK0_SB2_n15), .A(
        EK0_SB2_n333), .B(EK0_SB2_n334), .ZN(EK0_SB2_n329) );
  OAI211_X1 EK0_SB2_U223 ( .C1(EK0_SB2_n462), .C2(EK0_SB2_n69), .A(EK0_SB2_n78), .B(EK0_SB2_n66), .ZN(EK0_SB2_n330) );
  AOI21_X1 EK0_SB2_U222 ( .B1(EK0_SB2_n327), .B2(EK0_SB2_n142), .A(EK0_SB2_n77), .ZN(EK0_SB2_n457) );
  OAI21_X1 EK0_SB2_U221 ( .B1(EK0_SB2_n231), .B2(EK0_SB2_n116), .A(
        EK0_SB2_n135), .ZN(EK0_SB2_n352) );
  AOI21_X1 EK0_SB2_U220 ( .B1(EK0_SB2_n172), .B2(EK0_SB2_n453), .A(
        EK0_SB2_n168), .ZN(EK0_SB2_n351) );
  OAI211_X1 EK0_SB2_U219 ( .C1(EK0_SB2_n351), .C2(EK0_SB2_n45), .A(
        EK0_SB2_n352), .B(EK0_SB2_n353), .ZN(EK0_SB2_n343) );
  INV_X1 EK0_SB2_U218 ( .A(EK0_SB2_n159), .ZN(EK0_SB2_n14) );
  OAI21_X1 EK0_SB2_U217 ( .B1(EK0_SB2_n160), .B2(EK0_SB2_n161), .A(
        EK0_SB2_n133), .ZN(EK0_SB2_n158) );
  OAI211_X1 EK0_SB2_U216 ( .C1(EK0_SB2_n68), .C2(EK0_SB2_n33), .A(EK0_SB2_n158), .B(EK0_SB2_n14), .ZN(EK0_SB2_n150) );
  INV_X1 EK0_SB2_U215 ( .A(EK0_SB2_n121), .ZN(EK0_SB2_n76) );
  AOI21_X1 EK0_SB2_U214 ( .B1(EK0_SB2_n113), .B2(EK0_SB2_n114), .A(EK0_SB2_n78), .ZN(EK0_SB2_n112) );
  OAI21_X1 EK0_SB2_U213 ( .B1(EK0_SB2_n105), .B2(EK0_SB2_n171), .A(
        EK0_SB2_n172), .ZN(EK0_SB2_n170) );
  INV_X1 EK0_SB2_U212 ( .A(EK0_SB2_n102), .ZN(EK0_SB2_n37) );
  NAND2_X1 EK0_SB2_U211 ( .A1(EK0_SB2_n281), .A2(EK0_SB2_n110), .ZN(
        EK0_SB2_n115) );
  NOR2_X1 EK0_SB2_U210 ( .A1(EK0_SB2_n83), .A2(EK0_SB2_n231), .ZN(EK0_SB2_n250) );
  INV_X1 EK0_SB2_U209 ( .A(EK0_SB2_n148), .ZN(EK0_SB2_n39) );
  AOI22_X1 EK0_SB2_U208 ( .A1(EK0_SB2_n120), .A2(EK0_SB2_n117), .B1(
        EK0_SB2_n148), .B2(EK0_SB2_n149), .ZN(EK0_SB2_n147) );
  OAI211_X1 EK0_SB2_U207 ( .C1(EK0_SB2_n84), .C2(EK0_SB2_n145), .A(
        EK0_SB2_n146), .B(EK0_SB2_n147), .ZN(EK0_SB2_n127) );
  INV_X1 EK0_SB2_U206 ( .A(EK0_SB2_n110), .ZN(EK0_SB2_n56) );
  NOR2_X1 EK0_SB2_U205 ( .A1(EK0_SB2_n50), .A2(EK0_SB2_n55), .ZN(EK0_SB2_n125)
         );
  NOR2_X1 EK0_SB2_U204 ( .A1(EK0_SB2_n120), .A2(EK0_SB2_n121), .ZN(
        EK0_SB2_n101) );
  AOI221_X1 EK0_SB2_U203 ( .B1(EK0_SB2_n190), .B2(EK0_SB2_n187), .C1(
        EK0_SB2_n264), .C2(EK0_SB2_n126), .A(EK0_SB2_n283), .ZN(EK0_SB2_n272)
         );
  NOR4_X1 EK0_SB2_U202 ( .A1(EK0_SB2_n274), .A2(EK0_SB2_n275), .A3(
        EK0_SB2_n276), .A4(EK0_SB2_n242), .ZN(EK0_SB2_n273) );
  AOI221_X1 EK0_SB2_U201 ( .B1(EK0_SB2_n311), .B2(EK0_SB2_n36), .C1(
        EK0_SB2_n312), .C2(EK0_SB2_n236), .A(EK0_SB2_n313), .ZN(EK0_SB2_n270)
         );
  NAND4_X1 EK0_SB2_U200 ( .A1(EK0_SB2_n270), .A2(EK0_SB2_n271), .A3(
        EK0_SB2_n272), .A4(EK0_SB2_n273), .ZN(EK0_n282) );
  NAND2_X1 EK0_SB2_U199 ( .A1(EK0_SB2_n48), .A2(EK0_SB2_n60), .ZN(EK0_SB2_n420) );
  AOI22_X1 EK0_SB2_U198 ( .A1(EK0_SB2_n231), .A2(EK0_SB2_n420), .B1(
        EK0_SB2_n219), .B2(EK0_SB2_n297), .ZN(EK0_SB2_n419) );
  AOI22_X1 EK0_SB2_U197 ( .A1(EK0_SB2_n219), .A2(EK0_SB2_n126), .B1(
        EK0_SB2_n137), .B2(EK0_SB2_n136), .ZN(EK0_SB2_n303) );
  INV_X1 EK0_SB2_U196 ( .A(EK0_SB2_n221), .ZN(EK0_SB2_n44) );
  NAND2_X1 EK0_SB2_U195 ( .A1(EK0_SB2_n143), .A2(EK0_SB2_n408), .ZN(
        EK0_SB2_n267) );
  NOR2_X1 EK0_SB2_U194 ( .A1(EK0_SB2_n7), .A2(EK0_SB2_n47), .ZN(EK0_SB2_n244)
         );
  INV_X1 EK0_SB2_U193 ( .A(EK0_SB2_n460), .ZN(EK0_SB2_n453) );
  AOI211_X1 EK0_SB2_U192 ( .C1(EK0_SB2_n231), .C2(EK0_SB2_n455), .A(
        EK0_SB2_n456), .B(EK0_SB2_n457), .ZN(EK0_SB2_n428) );
  AOI221_X1 EK0_SB2_U191 ( .B1(EK0_SB2_n454), .B2(EK0_SB2_n324), .C1(
        EK0_SB2_n401), .C2(EK0_SB2_n149), .A(EK0_SB2_n458), .ZN(EK0_SB2_n427)
         );
  NAND4_X1 EK0_SB2_U190 ( .A1(EK0_SB2_n427), .A2(EK0_SB2_n428), .A3(
        EK0_SB2_n429), .A4(EK0_SB2_n430), .ZN(EK0_n278) );
  OAI22_X1 EK0_SB2_U189 ( .A1(EK0_SB2_n182), .A2(EK0_SB2_n76), .B1(EK0_SB2_n71), .B2(EK0_SB2_n29), .ZN(EK0_SB2_n262) );
  AOI21_X1 EK0_SB2_U188 ( .B1(EK0_SB2_n137), .B2(EK0_SB2_n462), .A(
        EK0_SB2_n126), .ZN(EK0_SB2_n215) );
  OAI22_X1 EK0_SB2_U187 ( .A1(EK0_SB2_n49), .A2(EK0_SB2_n74), .B1(EK0_SB2_n215), .B2(EK0_SB2_n80), .ZN(EK0_SB2_n214) );
  OAI22_X1 EK0_SB2_U186 ( .A1(EK0_SB2_n41), .A2(EK0_SB2_n56), .B1(EK0_SB2_n59), 
        .B2(EK0_SB2_n37), .ZN(EK0_SB2_n368) );
  AOI22_X1 EK0_SB2_U185 ( .A1(EK0_SB2_n36), .A2(EK0_SB2_n453), .B1(
        EK0_SB2_n202), .B2(EK0_SB2_n85), .ZN(EK0_SB2_n266) );
  OAI221_X1 EK0_SB2_U184 ( .B1(EK0_SB2_n453), .B2(EK0_SB2_n29), .C1(
        EK0_SB2_n462), .C2(EK0_SB2_n33), .A(EK0_SB2_n266), .ZN(EK0_SB2_n265)
         );
  OAI22_X1 EK0_SB2_U183 ( .A1(EK0_SB2_n55), .A2(EK0_SB2_n75), .B1(EK0_SB2_n56), 
        .B2(EK0_SB2_n73), .ZN(EK0_SB2_n374) );
  NOR3_X1 EK0_SB2_U182 ( .A1(EK0_SB2_n65), .A2(EK0_SB2_n461), .A3(EK0_SB2_n50), 
        .ZN(EK0_SB2_n375) );
  AOI21_X1 EK0_SB2_U181 ( .B1(EK0_SB2_n459), .B2(EK0_SB2_n367), .A(EK0_SB2_n51), .ZN(EK0_SB2_n376) );
  NOR3_X1 EK0_SB2_U180 ( .A1(EK0_SB2_n374), .A2(EK0_SB2_n375), .A3(
        EK0_SB2_n376), .ZN(EK0_SB2_n373) );
  INV_X1 EK0_SB2_U179 ( .A(EK0_SB2_n124), .ZN(EK0_SB2_n73) );
  NOR2_X1 EK0_SB2_U178 ( .A1(EK0_SB2_n68), .A2(EK0_SB2_n460), .ZN(EK0_SB2_n190) );
  NOR2_X1 EK0_SB2_U177 ( .A1(EK0_SB2_n141), .A2(EK0_SB2_n7), .ZN(EK0_SB2_n277)
         );
  INV_X1 EK0_SB2_U176 ( .A(EK0_SB2_n172), .ZN(EK0_SB2_n62) );
  AOI21_X1 EK0_SB2_U175 ( .B1(EK0_SB2_n70), .B2(EK0_SB2_n78), .A(EK0_SB2_n34), 
        .ZN(EK0_SB2_n320) );
  OAI21_X1 EK0_SB2_U174 ( .B1(EK0_SB2_n197), .B2(EK0_SB2_n327), .A(
        EK0_SB2_n328), .ZN(EK0_SB2_n318) );
  AOI211_X1 EK0_SB2_U173 ( .C1(EK0_SB2_n318), .C2(EK0_SB2_n462), .A(
        EK0_SB2_n319), .B(EK0_SB2_n320), .ZN(EK0_SB2_n317) );
  AOI21_X1 EK0_SB2_U172 ( .B1(EK0_SB2_n68), .B2(EK0_SB2_n76), .A(EK0_SB2_n6), 
        .ZN(EK0_SB2_n97) );
  NOR3_X1 EK0_SB2_U171 ( .A1(EK0_SB2_n85), .A2(EK0_SB2_n57), .A3(EK0_SB2_n37), 
        .ZN(EK0_SB2_n96) );
  NOR4_X1 EK0_SB2_U170 ( .A1(EK0_SB2_n94), .A2(EK0_SB2_n95), .A3(EK0_SB2_n96), 
        .A4(EK0_SB2_n97), .ZN(EK0_SB2_n93) );
  NOR2_X1 EK0_SB2_U169 ( .A1(EK0_SB2_n172), .A2(EK0_SB2_n312), .ZN(
        EK0_SB2_n197) );
  NOR2_X1 EK0_SB2_U168 ( .A1(EK0_SB2_n45), .A2(EK0_SB2_n7), .ZN(EK0_SB2_n161)
         );
  INV_X1 EK0_SB2_U167 ( .A(EK0_SB2_n126), .ZN(EK0_SB2_n60) );
  OAI221_X1 EK0_SB2_U166 ( .B1(EK0_SB2_n49), .B2(EK0_SB2_n78), .C1(EK0_SB2_n81), .C2(EK0_SB2_n60), .A(EK0_SB2_n369), .ZN(EK0_SB2_n361) );
  NOR2_X1 EK0_SB2_U165 ( .A1(EK0_SB2_n44), .A2(EK0_SB2_n7), .ZN(EK0_SB2_n217)
         );
  INV_X1 EK0_SB2_U164 ( .A(EK0_SB2_n256), .ZN(EK0_SB2_n46) );
  OAI221_X1 EK0_SB2_U163 ( .B1(EK0_SB2_n73), .B2(EK0_SB2_n54), .C1(EK0_SB2_n50), .C2(EK0_SB2_n79), .A(EK0_SB2_n341), .ZN(EK0_SB2_n335) );
  OAI21_X1 EK0_SB2_U162 ( .B1(EK0_SB2_n137), .B2(EK0_SB2_n171), .A(
        EK0_SB2_n219), .ZN(EK0_SB2_n407) );
  OAI221_X1 EK0_SB2_U161 ( .B1(EK0_SB2_n80), .B2(EK0_SB2_n141), .C1(
        EK0_SB2_n406), .C2(EK0_SB2_n84), .A(EK0_SB2_n407), .ZN(EK0_SB2_n405)
         );
  NOR2_X1 EK0_SB2_U160 ( .A1(EK0_SB2_n102), .A2(EK0_SB2_n221), .ZN(
        EK0_SB2_n220) );
  OAI221_X1 EK0_SB2_U159 ( .B1(EK0_SB2_n220), .B2(EK0_SB2_n62), .C1(
        EK0_SB2_n57), .C2(EK0_SB2_n35), .A(EK0_SB2_n8), .ZN(EK0_SB2_n218) );
  OAI21_X1 EK0_SB2_U158 ( .B1(EK0_SB2_n136), .B2(EK0_SB2_n462), .A(
        EK0_SB2_n259), .ZN(EK0_SB2_n412) );
  NOR2_X1 EK0_SB2_U157 ( .A1(EK0_SB2_n297), .A2(EK0_SB2_n135), .ZN(
        EK0_SB2_n411) );
  OAI221_X1 EK0_SB2_U156 ( .B1(EK0_SB2_n411), .B2(EK0_SB2_n73), .C1(
        EK0_SB2_n44), .C2(EK0_SB2_n61), .A(EK0_SB2_n412), .ZN(EK0_SB2_n410) );
  INV_X1 EK0_SB2_U155 ( .A(EK0_SB2_n298), .ZN(EK0_SB2_n51) );
  INV_X1 EK0_SB2_U154 ( .A(EK0_SB2_n259), .ZN(EK0_SB2_n54) );
  OAI221_X1 EK0_SB2_U153 ( .B1(EK0_SB2_n453), .B2(EK0_SB2_n6), .C1(EK0_SB2_n23), .C2(EK0_SB2_n88), .A(EK0_SB2_n146), .ZN(EK0_SB2_n325) );
  AOI221_X1 EK0_SB2_U152 ( .B1(EK0_SB2_n36), .B2(EK0_SB2_n231), .C1(
        EK0_SB2_n324), .C2(EK0_SB2_n460), .A(EK0_SB2_n325), .ZN(EK0_SB2_n322)
         );
  NAND2_X1 EK0_SB2_U151 ( .A1(EK0_SB2_n65), .A2(EK0_SB2_n72), .ZN(EK0_SB2_n299) );
  INV_X1 EK0_SB2_U150 ( .A(EK0_SB2_n300), .ZN(EK0_SB2_n52) );
  AOI221_X1 EK0_SB2_U149 ( .B1(EK0_SB2_n168), .B2(EK0_SB2_n297), .C1(
        EK0_SB2_n298), .C2(EK0_SB2_n299), .A(EK0_SB2_n52), .ZN(EK0_SB2_n293)
         );
  INV_X1 EK0_SB2_U148 ( .A(EK0_SB2_n243), .ZN(EK0_SB2_n25) );
  NOR4_X1 EK0_SB2_U147 ( .A1(EK0_SB2_n240), .A2(EK0_SB2_n25), .A3(EK0_SB2_n241), .A4(EK0_SB2_n242), .ZN(EK0_SB2_n239) );
  NOR2_X1 EK0_SB2_U146 ( .A1(EK0_SB2_n75), .A2(EK0_SB2_n462), .ZN(EK0_SB2_n173) );
  NOR3_X1 EK0_SB2_U145 ( .A1(EK0_SB2_n35), .A2(EK0_SB2_n47), .A3(EK0_SB2_n75), 
        .ZN(EK0_SB2_n241) );
  AOI21_X1 EK0_SB2_U144 ( .B1(EK0_SB2_n55), .B2(EK0_SB2_n307), .A(EK0_SB2_n86), 
        .ZN(EK0_SB2_n306) );
  NOR3_X1 EK0_SB2_U143 ( .A1(EK0_SB2_n75), .A2(EK0_SB2_n461), .A3(EK0_SB2_n49), 
        .ZN(EK0_SB2_n305) );
  AOI211_X1 EK0_SB2_U142 ( .C1(EK0_SB2_n269), .C2(EK0_SB2_n134), .A(
        EK0_SB2_n305), .B(EK0_SB2_n306), .ZN(EK0_SB2_n304) );
  OAI22_X1 EK0_SB2_U141 ( .A1(EK0_SB2_n462), .A2(EK0_SB2_n34), .B1(
        EK0_SB2_n460), .B2(EK0_SB2_n33), .ZN(EK0_SB2_n377) );
  AOI211_X1 EK0_SB2_U140 ( .C1(EK0_SB2_n339), .C2(EK0_SB2_n460), .A(
        EK0_SB2_n377), .B(EK0_SB2_n193), .ZN(EK0_SB2_n372) );
  NOR2_X1 EK0_SB2_U139 ( .A1(EK0_SB2_n56), .A2(EK0_SB2_n50), .ZN(EK0_SB2_n245)
         );
  INV_X1 EK0_SB2_U138 ( .A(EK0_SB2_n297), .ZN(EK0_SB2_n49) );
  OAI21_X1 EK0_SB2_U137 ( .B1(EK0_SB2_n57), .B2(EK0_SB2_n39), .A(EK0_SB2_n20), 
        .ZN(EK0_SB2_n399) );
  AOI21_X1 EK0_SB2_U136 ( .B1(EK0_SB2_n12), .B2(EK0_SB2_n312), .A(EK0_SB2_n132), .ZN(EK0_SB2_n397) );
  AOI21_X1 EK0_SB2_U135 ( .B1(EK0_SB2_n134), .B2(EK0_SB2_n399), .A(
        EK0_SB2_n400), .ZN(EK0_SB2_n398) );
  OAI221_X1 EK0_SB2_U134 ( .B1(EK0_SB2_n397), .B2(EK0_SB2_n462), .C1(
        EK0_SB2_n75), .C2(EK0_SB2_n8), .A(EK0_SB2_n398), .ZN(EK0_SB2_n392) );
  AOI21_X1 EK0_SB2_U133 ( .B1(EK0_SB2_n269), .B2(EK0_SB2_n281), .A(
        EK0_SB2_n282), .ZN(EK0_SB2_n279) );
  OAI21_X1 EK0_SB2_U132 ( .B1(EK0_SB2_n168), .B2(EK0_SB2_n116), .A(EK0_SB2_n31), .ZN(EK0_SB2_n280) );
  NAND2_X1 EK0_SB2_U131 ( .A1(EK0_SB2_n85), .A2(EK0_SB2_n70), .ZN(EK0_SB2_n278) );
  OAI221_X1 EK0_SB2_U130 ( .B1(EK0_SB2_n2), .B2(EK0_SB2_n278), .C1(
        EK0_SB2_n279), .C2(EK0_SB2_n84), .A(EK0_SB2_n280), .ZN(EK0_SB2_n274)
         );
  INV_X1 EK0_SB2_U129 ( .A(EK0_SB2_n123), .ZN(EK0_SB2_n68) );
  NOR2_X1 EK0_SB2_U128 ( .A1(EK0_SB2_n35), .A2(EK0_SB2_n44), .ZN(EK0_SB2_n202)
         );
  NOR2_X1 EK0_SB2_U127 ( .A1(EK0_SB2_n80), .A2(EK0_SB2_n462), .ZN(EK0_SB2_n116) );
  AOI221_X1 EK0_SB2_U126 ( .B1(EK0_SB2_n172), .B2(EK0_SB2_n231), .C1(
        EK0_SB2_n135), .C2(EK0_SB2_n288), .A(EK0_SB2_n405), .ZN(EK0_SB2_n404)
         );
  AOI221_X1 EK0_SB2_U125 ( .B1(EK0_SB2_n408), .B2(EK0_SB2_n409), .C1(
        EK0_SB2_n135), .C2(EK0_SB2_n231), .A(EK0_SB2_n410), .ZN(EK0_SB2_n403)
         );
  OAI222_X1 EK0_SB2_U124 ( .A1(EK0_SB2_n403), .A2(EK0_SB2_n7), .B1(
        EK0_SB2_n404), .B2(EK0_SB2_n30), .C1(EK0_SB2_n29), .C2(EK0_SB2_n69), 
        .ZN(EK0_SB2_n402) );
  INV_X1 EK0_SB2_U123 ( .A(EK0_SB2_n132), .ZN(EK0_SB2_n16) );
  AOI222_X1 EK0_SB2_U122 ( .A1(EK0_SB2_n133), .A2(EK0_SB2_n134), .B1(
        EK0_SB2_n135), .B2(EK0_SB2_n136), .C1(EK0_SB2_n137), .C2(EK0_SB2_n124), 
        .ZN(EK0_SB2_n131) );
  OAI222_X1 EK0_SB2_U121 ( .A1(EK0_SB2_n48), .A2(EK0_SB2_n130), .B1(
        EK0_SB2_n131), .B2(EK0_SB2_n7), .C1(EK0_SB2_n86), .C2(EK0_SB2_n16), 
        .ZN(EK0_SB2_n129) );
  AOI22_X1 EK0_SB2_U120 ( .A1(EK0_SB2_n157), .A2(EK0_SB2_n221), .B1(
        EK0_SB2_n136), .B2(EK0_SB2_n50), .ZN(EK0_SB2_n296) );
  OAI222_X1 EK0_SB2_U119 ( .A1(EK0_SB2_n49), .A2(EK0_SB2_n80), .B1(
        EK0_SB2_n461), .B2(EK0_SB2_n296), .C1(EK0_SB2_n55), .C2(EK0_SB2_n74), 
        .ZN(EK0_SB2_n295) );
  AOI221_X1 EK0_SB2_U118 ( .B1(EK0_SB2_n126), .B2(EK0_SB2_n287), .C1(
        EK0_SB2_n137), .C2(EK0_SB2_n144), .A(EK0_SB2_n295), .ZN(EK0_SB2_n294)
         );
  NOR2_X1 EK0_SB2_U117 ( .A1(EK0_SB2_n460), .A2(EK0_SB2_n70), .ZN(EK0_SB2_n312) );
  NOR4_X1 EK0_SB2_U116 ( .A1(EK0_SB2_n461), .A2(EK0_SB2_n41), .A3(EK0_SB2_n64), 
        .A4(EK0_SB2_n51), .ZN(EK0_SB2_n275) );
  NOR2_X1 EK0_SB2_U115 ( .A1(EK0_SB2_n50), .A2(EK0_SB2_n59), .ZN(EK0_SB2_n408)
         );
  NOR2_X1 EK0_SB2_U114 ( .A1(EK0_SB2_n51), .A2(EK0_SB2_n7), .ZN(EK0_SB2_n156)
         );
  NOR2_X1 EK0_SB2_U113 ( .A1(EK0_SB2_n51), .A2(EK0_SB2_n35), .ZN(EK0_SB2_n324)
         );
  NOR2_X1 EK0_SB2_U112 ( .A1(EK0_SB2_n41), .A2(EK0_SB2_n50), .ZN(EK0_SB2_n103)
         );
  NOR2_X1 EK0_SB2_U111 ( .A1(EK0_SB2_n83), .A2(EK0_SB2_n59), .ZN(EK0_SB2_n288)
         );
  OAI22_X1 EK0_SB2_U110 ( .A1(EK0_SB2_n73), .A2(EK0_SB2_n115), .B1(
        EK0_SB2_n435), .B2(EK0_SB2_n462), .ZN(EK0_SB2_n434) );
  OAI222_X1 EK0_SB2_U109 ( .A1(EK0_SB2_n76), .A2(EK0_SB2_n342), .B1(EK0_U9_Z_0), .B2(EK0_SB2_n447), .C1(EK0_SB2_n459), .C2(EK0_SB2_n238), .ZN(EK0_SB2_n432)
         );
  OAI222_X1 EK0_SB2_U108 ( .A1(EK0_SB2_n42), .A2(EK0_SB2_n30), .B1(EK0_SB2_n64), .B2(EK0_SB2_n146), .C1(EK0_SB2_n449), .C2(EK0_SB2_n79), .ZN(EK0_SB2_n431) );
  NOR4_X1 EK0_SB2_U107 ( .A1(EK0_SB2_n431), .A2(EK0_SB2_n432), .A3(
        EK0_SB2_n433), .A4(EK0_SB2_n434), .ZN(EK0_SB2_n430) );
  INV_X1 EK0_SB2_U106 ( .A(EK0_SB2_n120), .ZN(EK0_SB2_n75) );
  NOR2_X2 EK0_SB2_U105 ( .A1(EK0_SB2_n460), .A2(EK0_SB2_n462), .ZN(
        EK0_SB2_n134) );
  NOR3_X1 EK0_SB2_U104 ( .A1(EK0_SB2_n85), .A2(EK0_SB2_n59), .A3(EK0_SB2_n4), 
        .ZN(EK0_SB2_n242) );
  NOR2_X1 EK0_SB2_U103 ( .A1(EK0_SB2_n462), .A2(EK0_SB2_n83), .ZN(EK0_SB2_n149) );
  NOR2_X2 EK0_SB2_U102 ( .A1(EK0_SB2_n460), .A2(EK0_SB2_n461), .ZN(
        EK0_SB2_n231) );
  NOR2_X1 EK0_SB2_U101 ( .A1(EK0_SB2_n460), .A2(EK0_SB2_n83), .ZN(EK0_SB2_n144) );
  NOR2_X1 EK0_SB2_U100 ( .A1(EK0_SB2_n462), .A2(EK0_SB2_n453), .ZN(
        EK0_SB2_n105) );
  NOR2_X1 EK0_SB2_U99 ( .A1(EK0_SB2_n50), .A2(EK0_SB2_n70), .ZN(EK0_SB2_n137)
         );
  NOR2_X1 EK0_SB2_U98 ( .A1(EK0_SB2_n83), .A2(EK0_SB2_n453), .ZN(EK0_SB2_n136)
         );
  INV_X1 EK0_SB2_U97 ( .A(EK0_SB2_n190), .ZN(EK0_SB2_n67) );
  INV_X1 EK0_SB2_U96 ( .A(EK0_SB2_n114), .ZN(EK0_SB2_n40) );
  AND2_X1 EK0_SB2_U95 ( .A1(EK0_SB2_n149), .A2(EK0_SB2_n244), .ZN(EK0_SB2_n360) );
  INV_X1 EK0_SB2_U94 ( .A(EK0_SB2_n396), .ZN(EK0_SB2_n27) );
  NAND2_X1 EK0_SB2_U93 ( .A1(EK0_SB2_n23), .A2(EK0_SB2_n39), .ZN(EK0_SB2_n379)
         );
  OR3_X1 EK0_SB2_U92 ( .A1(EK0_SB2_n49), .A2(EK0_SB2_n101), .A3(EK0_SB2_n23), 
        .ZN(EK0_SB2_n100) );
  INV_X1 EK0_SB2_U91 ( .A(EK0_SB2_n413), .ZN(EK0_SB2_n63) );
  INV_X1 EK0_SB2_U90 ( .A(EK0_SB2_n217), .ZN(EK0_SB2_n6) );
  INV_X1 EK0_SB2_U89 ( .A(EK0_SB2_n277), .ZN(EK0_SB2_n4) );
  INV_X1 EK0_SB2_U88 ( .A(EK0_SB2_n342), .ZN(EK0_SB2_n24) );
  INV_X1 EK0_SB2_U87 ( .A(EK0_SB2_n125), .ZN(EK0_SB2_n47) );
  NAND2_X1 EK0_SB2_U86 ( .A1(EK0_SB2_n39), .A2(EK0_SB2_n11), .ZN(EK0_SB2_n187)
         );
  NAND2_X1 EK0_SB2_U85 ( .A1(EK0_SB2_n134), .A2(EK0_SB2_n244), .ZN(
        EK0_SB2_n199) );
  NAND2_X1 EK0_SB2_U84 ( .A1(EK0_SB2_n77), .A2(EK0_SB2_n88), .ZN(EK0_SB2_n192)
         );
  INV_X1 EK0_SB2_U83 ( .A(EK0_SB2_n116), .ZN(EK0_SB2_n79) );
  INV_X1 EK0_SB2_U82 ( .A(EK0_SB2_n156), .ZN(EK0_SB2_n5) );
  INV_X1 EK0_SB2_U81 ( .A(EK0_SB2_n327), .ZN(EK0_SB2_n12) );
  INV_X1 EK0_SB2_U80 ( .A(EK0_SB2_n288), .ZN(EK0_SB2_n57) );
  NAND2_X1 EK0_SB2_U79 ( .A1(EK0_SB2_n77), .A2(EK0_SB2_n84), .ZN(EK0_SB2_n167)
         );
  INV_X1 EK0_SB2_U78 ( .A(EK0_SB2_n103), .ZN(EK0_SB2_n38) );
  INV_X1 EK0_SB2_U77 ( .A(EK0_SB2_n202), .ZN(EK0_SB2_n34) );
  INV_X1 EK0_SB2_U76 ( .A(EK0_SB2_n324), .ZN(EK0_SB2_n33) );
  OAI21_X1 EK0_SB2_U75 ( .B1(EK0_SB2_n459), .B2(EK0_SB2_n68), .A(EK0_SB2_n64), 
        .ZN(EK0_SB2_n444) );
  OAI21_X1 EK0_SB2_U74 ( .B1(EK0_SB2_n9), .B2(EK0_SB2_n54), .A(EK0_SB2_n18), 
        .ZN(EK0_SB2_n260) );
  OAI21_X1 EK0_SB2_U73 ( .B1(EK0_SB2_n66), .B2(EK0_SB2_n18), .A(EK0_SB2_n115), 
        .ZN(EK0_SB2_n109) );
  INV_X1 EK0_SB2_U72 ( .A(EK0_SB2_n173), .ZN(EK0_SB2_n74) );
  INV_X1 EK0_SB2_U71 ( .A(EK0_SB2_n137), .ZN(EK0_SB2_n48) );
  INV_X1 EK0_SB2_U70 ( .A(EK0_SB2_n185), .ZN(EK0_SB2_n55) );
  AOI21_X1 EK0_SB2_U69 ( .B1(EK0_SB2_n88), .B2(EK0_SB2_n80), .A(EK0_SB2_n115), 
        .ZN(EK0_SB2_n366) );
  AOI21_X1 EK0_SB2_U68 ( .B1(EK0_SB2_n82), .B2(EK0_SB2_n78), .A(EK0_SB2_n23), 
        .ZN(EK0_SB2_n119) );
  INV_X1 EK0_SB2_U67 ( .A(EK0_SB2_n231), .ZN(EK0_SB2_n86) );
  NOR2_X1 EK0_SB2_U66 ( .A1(EK0_SB2_n60), .A2(EK0_SB2_n9), .ZN(EK0_SB2_n401)
         );
  INV_X1 EK0_SB2_U65 ( .A(EK0_SB2_n267), .ZN(EK0_SB2_n31) );
  INV_X1 EK0_SB2_U64 ( .A(EK0_SB2_n311), .ZN(EK0_SB2_n69) );
  NOR2_X1 EK0_SB2_U63 ( .A1(EK0_SB2_n71), .A2(EK0_SB2_n15), .ZN(EK0_SB2_n240)
         );
  NOR2_X1 EK0_SB2_U62 ( .A1(EK0_SB2_n62), .A2(EK0_SB2_n453), .ZN(EK0_SB2_n445)
         );
  INV_X1 EK0_SB2_U61 ( .A(EK0_SB2_n312), .ZN(EK0_SB2_n65) );
  NOR2_X1 EK0_SB2_U60 ( .A1(EK0_SB2_n51), .A2(EK0_SB2_n30), .ZN(EK0_SB2_n381)
         );
  INV_X1 EK0_SB2_U59 ( .A(EK0_SB2_n161), .ZN(EK0_SB2_n2) );
  INV_X1 EK0_SB2_U58 ( .A(EK0_SB2_n157), .ZN(EK0_SB2_n66) );
  INV_X1 EK0_SB2_U57 ( .A(EK0_SB2_n134), .ZN(EK0_SB2_n85) );
  INV_X1 EK0_SB2_U56 ( .A(EK0_SB2_n144), .ZN(EK0_SB2_n82) );
  OAI22_X1 EK0_SB2_U55 ( .A1(EK0_SB2_n38), .A2(EK0_SB2_n80), .B1(EK0_SB2_n39), 
        .B2(EK0_SB2_n81), .ZN(EK0_SB2_n111) );
  OAI22_X1 EK0_SB2_U54 ( .A1(EK0_SB2_n55), .A2(EK0_SB2_n79), .B1(EK0_SB2_n459), 
        .B2(EK0_SB2_n54), .ZN(EK0_SB2_n261) );
  AOI21_X1 EK0_SB2_U53 ( .B1(EK0_SB2_n45), .B2(EK0_SB2_n68), .A(EK0_SB2_n130), 
        .ZN(EK0_SB2_n228) );
  OAI22_X1 EK0_SB2_U52 ( .A1(EK0_SB2_n56), .A2(EK0_SB2_n75), .B1(EK0_SB2_n81), 
        .B2(EK0_SB2_n48), .ZN(EK0_SB2_n446) );
  OAI22_X1 EK0_SB2_U51 ( .A1(EK0_SB2_n82), .A2(EK0_SB2_n18), .B1(EK0_SB2_n461), 
        .B2(EK0_SB2_n267), .ZN(EK0_SB2_n383) );
  NOR2_X1 EK0_SB2_U50 ( .A1(EK0_SB2_n18), .A2(EK0_SB2_n461), .ZN(EK0_SB2_n193)
         );
  NOR2_X1 EK0_SB2_U49 ( .A1(EK0_SB2_n45), .A2(EK0_SB2_n23), .ZN(EK0_SB2_n339)
         );
  NOR2_X1 EK0_SB2_U48 ( .A1(EK0_SB2_n141), .A2(EK0_SB2_n23), .ZN(EK0_SB2_n350)
         );
  NOR2_X1 EK0_SB2_U47 ( .A1(EK0_SB2_n60), .A2(EK0_SB2_n23), .ZN(EK0_SB2_n282)
         );
  NOR2_X1 EK0_SB2_U46 ( .A1(EK0_SB2_n82), .A2(EK0_SB2_n461), .ZN(EK0_SB2_n207)
         );
  NOR2_X1 EK0_SB2_U45 ( .A1(EK0_SB2_n15), .A2(EK0_SB2_n68), .ZN(EK0_SB2_n159)
         );
  OAI221_X1 EK0_SB2_U44 ( .B1(EK0_SB2_n49), .B2(EK0_SB2_n75), .C1(EK0_SB2_n86), 
        .C2(EK0_SB2_n64), .A(EK0_SB2_n300), .ZN(EK0_SB2_n362) );
  NOR2_X1 EK0_SB2_U43 ( .A1(EK0_SB2_n43), .A2(EK0_SB2_n23), .ZN(EK0_SB2_n188)
         );
  INV_X1 EK0_SB2_U42 ( .A(EK0_SB2_n136), .ZN(EK0_SB2_n80) );
  OAI222_X1 EK0_SB2_U41 ( .A1(EK0_SB2_n68), .A2(EK0_SB2_n33), .B1(EK0_SB2_n78), 
        .B2(EK0_SB2_n15), .C1(EK0_SB2_n77), .C2(EK0_SB2_n19), .ZN(EK0_SB2_n313) );
  NOR3_X1 EK0_SB2_U40 ( .A1(EK0_SB2_n72), .A2(EK0_SB2_n55), .A3(EK0_SB2_n39), 
        .ZN(EK0_SB2_n394) );
  INV_X1 EK0_SB2_U39 ( .A(EK0_SB2_n149), .ZN(EK0_SB2_n78) );
  INV_X1 EK0_SB2_U38 ( .A(EK0_SB2_n105), .ZN(EK0_SB2_n84) );
  NOR2_X1 EK0_SB2_U37 ( .A1(EK0_SB2_n51), .A2(EK0_SB2_n23), .ZN(EK0_SB2_n162)
         );
  NOR2_X1 EK0_SB2_U36 ( .A1(EK0_SB2_n44), .A2(EK0_SB2_n23), .ZN(EK0_SB2_n236)
         );
  AOI22_X1 EK0_SB2_U35 ( .A1(EK0_SB2_n157), .A2(EK0_SB2_n453), .B1(
        EK0_SB2_n144), .B2(EK0_SB2_n461), .ZN(EK0_SB2_n216) );
  OAI222_X1 EK0_SB2_U34 ( .A1(EK0_SB2_n48), .A2(EK0_SB2_n75), .B1(EK0_SB2_n216), .B2(EK0_SB2_n45), .C1(EK0_SB2_n459), .C2(EK0_SB2_n55), .ZN(EK0_SB2_n211) );
  NOR2_X1 EK0_SB2_U33 ( .A1(EK0_SB2_n30), .A2(EK0_SB2_n44), .ZN(EK0_SB2_n160)
         );
  NOR2_X1 EK0_SB2_U32 ( .A1(EK0_U9_Z_0), .A2(EK0_SB2_n453), .ZN(EK0_SB2_n287)
         );
  NOR2_X1 EK0_SB2_U31 ( .A1(EK0_SB2_n73), .A2(EK0_SB2_n461), .ZN(EK0_SB2_n168)
         );
  INV_X1 EK0_SB2_U30 ( .A(EK0_SB2_n381), .ZN(EK0_SB2_n28) );
  INV_X1 EK0_SB2_U29 ( .A(EK0_SB2_n193), .ZN(EK0_SB2_n17) );
  INV_X1 EK0_SB2_U28 ( .A(EK0_SB2_n445), .ZN(EK0_SB2_n61) );
  INV_X1 EK0_SB2_U27 ( .A(EK0_SB2_n401), .ZN(EK0_SB2_n8) );
  INV_X1 EK0_SB2_U26 ( .A(EK0_SB2_n350), .ZN(EK0_SB2_n21) );
  INV_X1 EK0_SB2_U25 ( .A(EK0_SB2_n162), .ZN(EK0_SB2_n20) );
  INV_X1 EK0_SB2_U24 ( .A(EK0_SB2_n188), .ZN(EK0_SB2_n19) );
  INV_X1 EK0_SB2_U23 ( .A(EK0_SB2_n160), .ZN(EK0_SB2_n29) );
  INV_X1 EK0_SB2_U22 ( .A(EK0_SB2_n236), .ZN(EK0_SB2_n18) );
  INV_X1 EK0_SB2_U21 ( .A(EK0_SB2_n168), .ZN(EK0_SB2_n72) );
  AOI21_X1 EK0_SB2_U20 ( .B1(EK0_SB2_n65), .B2(EK0_SB2_n61), .A(EK0_SB2_n2), 
        .ZN(EK0_SB2_n456) );
  AOI21_X1 EK0_SB2_U19 ( .B1(EK0_SB2_n85), .B2(EK0_SB2_n63), .A(EK0_SB2_n34), 
        .ZN(EK0_SB2_n458) );
  INV_X1 EK0_SB2_U18 ( .A(EK0_SB2_n207), .ZN(EK0_SB2_n81) );
  INV_X1 EK0_SB2_U17 ( .A(EK0_SB2_n339), .ZN(EK0_SB2_n15) );
  INV_X1 EK0_SB2_U16 ( .A(EK0_SB2_n287), .ZN(EK0_SB2_n88) );
  BUF_X2 EK0_SB2_U15 ( .A(EK0_U9_Z_2), .Z(EK0_SB2_n89) );
  INV_X1 EK0_SB2_U14 ( .A(EK0_U9_Z_3), .ZN(EK0_SB2_n70) );
  NOR2_X1 EK0_SB2_U13 ( .A1(EK0_SB2_n70), .A2(EK0_U9_Z_4), .ZN(EK0_SB2_n126)
         );
  NOR2_X1 EK0_SB2_U12 ( .A1(EK0_SB2_n70), .A2(EK0_SB2_n452), .ZN(EK0_SB2_n135)
         );
  NOR2_X1 EK0_SB2_U11 ( .A1(EK0_SB2_n32), .A2(EK0_n569), .ZN(EK0_SB2_n143) );
  BUF_X2 EK0_SB2_U10 ( .A(EK0_U9_Z_5), .Z(EK0_SB2_n452) );
  INV_X1 EK0_SB2_U9 ( .A(EK0_SB2_n163), .ZN(EK0_SB2_n35) );
  INV_X1 EK0_SB2_U8 ( .A(EK0_SB2_n133), .ZN(EK0_SB2_n64) );
  INV_X1 EK0_SB2_U7 ( .A(EK0_n286), .ZN(EK0_SB2_n32) );
  INV_X1 EK0_SB2_U6 ( .A(EK0_SB2_n143), .ZN(EK0_SB2_n30) );
  NOR2_X1 EK0_SB2_U5 ( .A1(EK0_SB2_n50), .A2(EK0_U9_Z_4), .ZN(EK0_SB2_n171) );
  NOR2_X1 EK0_SB2_U4 ( .A1(EK0_SB2_n32), .A2(EK0_SB2_n41), .ZN(EK0_SB2_n246)
         );
  NOR2_X1 EK0_SB2_U3 ( .A1(EK0_SB2_n41), .A2(EK0_n286), .ZN(EK0_SB2_n163) );
  INV_X2 EK0_SB2_U2 ( .A(EK0_U9_Z_4), .ZN(EK0_SB2_n59) );
  INV_X2 EK0_SB2_U1 ( .A(EK0_SB2_n246), .ZN(EK0_SB2_n23) );
  NAND3_X1 EK0_SB2_U464 ( .A1(EK0_SB2_n143), .A2(EK0_SB2_n245), .A3(
        EK0_SB2_n121), .ZN(EK0_SB2_n396) );
  OAI33_X1 EK0_SB2_U463 ( .A1(EK0_SB2_n75), .A2(EK0_SB2_n55), .A3(EK0_SB2_n7), 
        .B1(EK0_SB2_n60), .B2(EK0_SB2_n83), .B3(EK0_SB2_n39), .ZN(EK0_SB2_n448) );
  NAND3_X1 EK0_SB2_U462 ( .A1(EK0_SB2_n408), .A2(EK0_SB2_n213), .A3(
        EK0_SB2_n157), .ZN(EK0_SB2_n238) );
  OAI33_X1 EK0_SB2_U461 ( .A1(EK0_SB2_n85), .A2(EK0_n286), .A3(EK0_SB2_n89), 
        .B1(EK0_SB2_n443), .B2(EK0_SB2_n59), .B3(EK0_SB2_n84), .ZN(
        EK0_SB2_n442) );
  NAND3_X1 EK0_SB2_U459 ( .A1(EK0_SB2_n134), .A2(EK0_SB2_n89), .A3(
        EK0_SB2_n117), .ZN(EK0_SB2_n421) );
  NAND4_X1 EK0_SB2_U458 ( .A1(EK0_SB2_n172), .A2(EK0_SB2_n287), .A3(
        EK0_SB2_n148), .A4(EK0_n286), .ZN(EK0_SB2_n422) );
  NAND3_X1 EK0_SB2_U457 ( .A1(EK0_SB2_n102), .A2(EK0_SB2_n83), .A3(
        EK0_SB2_n231), .ZN(EK0_SB2_n423) );
  NAND3_X1 EK0_SB2_U456 ( .A1(EK0_SB2_n421), .A2(EK0_SB2_n422), .A3(
        EK0_SB2_n423), .ZN(EK0_SB2_n417) );
  NAND3_X1 EK0_SB2_U455 ( .A1(EK0_SB2_n69), .A2(EK0_SB2_n77), .A3(EK0_SB2_n367), .ZN(EK0_SB2_n409) );
  OAI33_X1 EK0_SB2_U454 ( .A1(EK0_SB2_n86), .A2(EK0_SB2_n57), .A3(EK0_SB2_n9), 
        .B1(EK0_SB2_n15), .B2(EK0_SB2_n70), .B3(EK0_SB2_n88), .ZN(EK0_SB2_n400) );
  NAND3_X1 EK0_SB2_U453 ( .A1(EK0_SB2_n244), .A2(EK0_SB2_n462), .A3(
        EK0_SB2_n89), .ZN(EK0_SB2_n99) );
  NAND3_X1 EK0_SB2_U452 ( .A1(EK0_SB2_n245), .A2(EK0_SB2_n246), .A3(
        EK0_SB2_n136), .ZN(EK0_SB2_n243) );
  NAND3_X1 EK0_SB2_U451 ( .A1(EK0_SB2_n99), .A2(EK0_SB2_n396), .A3(
        EK0_SB2_n243), .ZN(EK0_SB2_n393) );
  OAI33_X1 EK0_SB2_U450 ( .A1(EK0_SB2_n81), .A2(EK0_SB2_n49), .A3(EK0_SB2_n23), 
        .B1(EK0_SB2_n84), .B2(EK0_n286), .B3(EK0_SB2_n47), .ZN(EK0_SB2_n395)
         );
  NAND3_X1 EK0_SB2_U448 ( .A1(EK0_SB2_n171), .A2(EK0_SB2_n312), .A3(
        EK0_SB2_n219), .ZN(EK0_SB2_n369) );
  NAND3_X1 EK0_SB2_U447 ( .A1(EK0_SB2_n231), .A2(EK0_SB2_n59), .A3(
        EK0_SB2_n206), .ZN(EK0_SB2_n333) );
  OAI33_X1 EK0_SB2_U446 ( .A1(EK0_SB2_n54), .A2(EK0_SB2_n83), .A3(EK0_SB2_n11), 
        .B1(EK0_SB2_n37), .B2(EK0_SB2_n459), .B3(EK0_SB2_n230), .ZN(
        EK0_SB2_n358) );
  NAND3_X1 EK0_SB2_U444 ( .A1(EK0_SB2_n83), .A2(EK0_SB2_n41), .A3(EK0_SB2_n206), .ZN(EK0_SB2_n349) );
  NAND4_X1 EK0_SB2_U443 ( .A1(EK0_SB2_n349), .A2(EK0_SB2_n19), .A3(
        EK0_SB2_n115), .A4(EK0_SB2_n267), .ZN(EK0_SB2_n346) );
  NAND3_X1 EK0_SB2_U442 ( .A1(EK0_SB2_n461), .A2(EK0_U9_Z_3), .A3(EK0_SB2_n171), .ZN(EK0_SB2_n256) );
  NAND3_X1 EK0_SB2_U441 ( .A1(EK0_SB2_n157), .A2(EK0_SB2_n59), .A3(
        EK0_SB2_n206), .ZN(EK0_SB2_n328) );
  NAND3_X1 EK0_SB2_U440 ( .A1(EK0_SB2_n172), .A2(EK0_SB2_n461), .A3(
        EK0_SB2_n31), .ZN(EK0_SB2_n323) );
  NAND4_X1 EK0_SB2_U439 ( .A1(EK0_SB2_n314), .A2(EK0_SB2_n315), .A3(
        EK0_SB2_n316), .A4(EK0_SB2_n317), .ZN(EK0_n281) );
  NAND3_X1 EK0_SB2_U437 ( .A1(EK0_SB2_n231), .A2(EK0_SB2_n70), .A3(
        EK0_SB2_n171), .ZN(EK0_SB2_n255) );
  NAND3_X1 EK0_SB2_U436 ( .A1(EK0_SB2_n461), .A2(EK0_SB2_n59), .A3(
        EK0_SB2_n123), .ZN(EK0_SB2_n257) );
  NAND4_X1 EK0_SB2_U435 ( .A1(EK0_SB2_n255), .A2(EK0_SB2_n256), .A3(
        EK0_SB2_n257), .A4(EK0_SB2_n258), .ZN(EK0_SB2_n247) );
  OAI33_X1 EK0_SB2_U434 ( .A1(EK0_SB2_n51), .A2(EK0_n286), .A3(EK0_SB2_n66), 
        .B1(EK0_SB2_n9), .B2(EK0_SB2_n55), .B3(EK0_SB2_n83), .ZN(EK0_SB2_n254)
         );
  NAND3_X1 EK0_SB2_U433 ( .A1(EK0_SB2_n245), .A2(EK0_SB2_n246), .A3(
        EK0_SB2_n149), .ZN(EK0_SB2_n198) );
  NAND4_X1 EK0_SB2_U432 ( .A1(EK0_SB2_n198), .A2(EK0_SB2_n199), .A3(
        EK0_SB2_n238), .A4(EK0_SB2_n239), .ZN(EK0_SB2_n226) );
  OAI33_X1 EK0_SB2_U431 ( .A1(EK0_SB2_n74), .A2(EK0_SB2_n43), .A3(EK0_SB2_n30), 
        .B1(EK0_SB2_n86), .B2(EK0_SB2_n230), .B3(EK0_SB2_n9), .ZN(EK0_SB2_n229) );
  NAND4_X1 EK0_SB2_U430 ( .A1(EK0_SB2_n222), .A2(EK0_SB2_n223), .A3(
        EK0_SB2_n224), .A4(EK0_SB2_n225), .ZN(EK0_n283) );
  NAND3_X1 EK0_SB2_U429 ( .A1(EK0_SB2_n68), .A2(EK0_SB2_n75), .A3(EK0_SB2_n84), 
        .ZN(EK0_SB2_n212) );
  OAI33_X1 EK0_SB2_U428 ( .A1(EK0_SB2_n37), .A2(EK0_SB2_n461), .A3(EK0_SB2_n83), .B1(EK0_SB2_n210), .B2(EK0_SB2_n78), .B3(EK0_SB2_n11), .ZN(EK0_SB2_n209) );
  NAND3_X1 EK0_SB2_U427 ( .A1(EK0_U9_Z_4), .A2(EK0_SB2_n201), .A3(EK0_n286), 
        .ZN(EK0_SB2_n200) );
  NAND3_X1 EK0_SB2_U426 ( .A1(EK0_SB2_n198), .A2(EK0_SB2_n199), .A3(
        EK0_SB2_n200), .ZN(EK0_SB2_n178) );
  NAND4_X1 EK0_SB2_U425 ( .A1(EK0_SB2_n174), .A2(EK0_SB2_n175), .A3(
        EK0_SB2_n176), .A4(EK0_SB2_n177), .ZN(EK0_n284) );
  NAND3_X1 EK0_SB2_U424 ( .A1(EK0_n286), .A2(EK0_SB2_n59), .A3(EK0_SB2_n120), 
        .ZN(EK0_SB2_n153) );
  NAND3_X1 EK0_SB2_U423 ( .A1(EK0_SB2_n152), .A2(EK0_SB2_n153), .A3(
        EK0_SB2_n154), .ZN(EK0_SB2_n151) );
  NAND3_X1 EK0_SB2_U422 ( .A1(EK0_n569), .A2(EK0_SB2_n59), .A3(EK0_SB2_n144), 
        .ZN(EK0_SB2_n138) );
  NAND3_X1 EK0_SB2_U421 ( .A1(EK0_SB2_n98), .A2(EK0_SB2_n99), .A3(EK0_SB2_n100), .ZN(EK0_SB2_n95) );
  NAND4_X1 EK0_SB2_U420 ( .A1(EK0_SB2_n90), .A2(EK0_SB2_n91), .A3(EK0_SB2_n92), 
        .A4(EK0_SB2_n93), .ZN(EK0_n285) );
  NOR2_X2 EK0_SB2_U313 ( .A1(EK0_SB2_n59), .A2(EK0_SB2_n70), .ZN(EK0_SB2_n185)
         );
  NOR2_X2 EK0_SB2_U264 ( .A1(EK0_SB2_n83), .A2(EK0_SB2_n70), .ZN(EK0_SB2_n157)
         );
  NOR2_X2 EK0_SB2_U263 ( .A1(EK0_SB2_n459), .A2(EK0_SB2_n89), .ZN(EK0_SB2_n120) );
endmodule

