
module mix_column ( data_in, data_out, rst, clk );
  input [127:0] data_in;
  output [127:0] data_out;
  input rst, clk;
  wire   n790, n792, n796, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;

  XOR2_X1 U38 ( .A(n802), .B(n803), .Z(data_out[9]) );
  XOR2_X1 U39 ( .A(n804), .B(n805), .Z(n803) );
  XOR2_X1 U40 ( .A(data_in[17]), .B(n806), .Z(n802) );
  XOR2_X1 U41 ( .A(n807), .B(n808), .Z(data_out[99]) );
  XOR2_X1 U42 ( .A(data_in[115]), .B(data_in[123]), .Z(n807) );
  XOR2_X1 U43 ( .A(n811), .B(n812), .Z(data_out[98]) );
  XOR2_X1 U44 ( .A(data_in[106]), .B(n813), .Z(n812) );
  XOR2_X1 U45 ( .A(data_in[97]), .B(data_in[105]), .Z(n811) );
  XOR2_X1 U46 ( .A(n814), .B(n815), .Z(data_out[97]) );
  XOR2_X1 U47 ( .A(n816), .B(n817), .Z(n815) );
  XOR2_X1 U48 ( .A(data_in[121]), .B(n818), .Z(n814) );
  XOR2_X1 U49 ( .A(n819), .B(n820), .Z(data_out[96]) );
  XOR2_X1 U50 ( .A(data_in[104]), .B(n821), .Z(n820) );
  XOR2_X1 U51 ( .A(n822), .B(n823), .Z(data_out[95]) );
  XOR2_X1 U52 ( .A(data_in[87]), .B(n824), .Z(n823) );
  XOR2_X1 U53 ( .A(n825), .B(n826), .Z(data_out[94]) );
  XOR2_X1 U54 ( .A(data_in[70]), .B(n827), .Z(n826) );
  XOR2_X1 U55 ( .A(n828), .B(n829), .Z(data_out[93]) );
  XOR2_X1 U56 ( .A(data_in[69]), .B(n830), .Z(n829) );
  XOR2_X1 U57 ( .A(n831), .B(n832), .Z(data_out[92]) );
  XOR2_X1 U58 ( .A(n833), .B(n834), .Z(n832) );
  XOR2_X1 U59 ( .A(data_in[68]), .B(n835), .Z(n831) );
  XOR2_X1 U62 ( .A(n840), .B(n841), .Z(data_out[90]) );
  XOR2_X1 U63 ( .A(data_in[82]), .B(n842), .Z(n841) );
  XOR2_X1 U64 ( .A(n843), .B(n844), .Z(data_out[8]) );
  XOR2_X1 U65 ( .A(data_in[0]), .B(n845), .Z(n844) );
  XOR2_X1 U66 ( .A(data_in[23]), .B(data_in[15]), .Z(n843) );
  XOR2_X1 U67 ( .A(n846), .B(n847), .Z(data_out[89]) );
  XOR2_X1 U68 ( .A(n848), .B(n849), .Z(n847) );
  XOR2_X1 U69 ( .A(data_in[65]), .B(n850), .Z(n846) );
  XOR2_X1 U70 ( .A(n851), .B(n852), .Z(data_out[88]) );
  XOR2_X1 U71 ( .A(data_in[80]), .B(n853), .Z(n852) );
  XOR2_X1 U72 ( .A(data_in[95]), .B(data_in[71]), .Z(n851) );
  XOR2_X1 U73 ( .A(n854), .B(n855), .Z(data_out[87]) );
  XOR2_X1 U74 ( .A(data_in[86]), .B(n822), .Z(n855) );
  XOR2_X1 U75 ( .A(data_in[95]), .B(data_in[94]), .Z(n854) );
  XOR2_X1 U76 ( .A(n856), .B(n857), .Z(data_out[86]) );
  XOR2_X1 U77 ( .A(data_in[78]), .B(n824), .Z(n857) );
  XOR2_X1 U78 ( .A(data_in[93]), .B(data_in[85]), .Z(n856) );
  XOR2_X1 U79 ( .A(n858), .B(n859), .Z(data_out[85]) );
  XOR2_X1 U80 ( .A(data_in[77]), .B(n827), .Z(n859) );
  XOR2_X1 U81 ( .A(data_in[92]), .B(data_in[84]), .Z(n858) );
  XOR2_X1 U82 ( .A(n860), .B(n861), .Z(data_out[84]) );
  XOR2_X1 U83 ( .A(n835), .B(n862), .Z(n861) );
  XOR2_X1 U84 ( .A(data_in[91]), .B(data_in[95]), .Z(n835) );
  XOR2_X1 U85 ( .A(data_in[76]), .B(n830), .Z(n860) );
  XOR2_X1 U86 ( .A(n863), .B(n864), .Z(data_out[83]) );
  XOR2_X1 U87 ( .A(data_in[90]), .B(data_in[95]), .Z(n837) );
  XOR2_X1 U88 ( .A(n866), .B(n867), .Z(data_out[82]) );
  XOR2_X1 U89 ( .A(data_in[90]), .B(n842), .Z(n867) );
  XOR2_X1 U90 ( .A(data_in[74]), .B(data_in[66]), .Z(n842) );
  XOR2_X1 U91 ( .A(data_in[89]), .B(data_in[81]), .Z(n866) );
  XOR2_X1 U92 ( .A(n868), .B(n869), .Z(data_out[81]) );
  XOR2_X1 U93 ( .A(n850), .B(n870), .Z(n869) );
  XOR2_X1 U94 ( .A(data_in[88]), .B(data_in[95]), .Z(n850) );
  XOR2_X1 U95 ( .A(data_in[73]), .B(n840), .Z(n868) );
  XOR2_X1 U96 ( .A(n871), .B(n872), .Z(data_out[80]) );
  XOR2_X1 U97 ( .A(data_in[88]), .B(n853), .Z(n872) );
  XOR2_X1 U98 ( .A(data_in[72]), .B(data_in[64]), .Z(n853) );
  XOR2_X1 U99 ( .A(n873), .B(n874), .Z(data_out[7]) );
  XOR2_X1 U100 ( .A(data_in[14]), .B(n875), .Z(n874) );
  XOR2_X1 U101 ( .A(data_in[6]), .B(data_in[15]), .Z(n873) );
  XOR2_X1 U102 ( .A(n871), .B(n876), .Z(data_out[79]) );
  XOR2_X1 U103 ( .A(data_in[71]), .B(n825), .Z(n876) );
  XOR2_X1 U104 ( .A(n828), .B(n877), .Z(data_out[78]) );
  XOR2_X1 U105 ( .A(data_in[86]), .B(n824), .Z(n877) );
  XOR2_X1 U106 ( .A(data_in[70]), .B(data_in[94]), .Z(n824) );
  XOR2_X1 U107 ( .A(n833), .B(n878), .Z(data_out[77]) );
  XOR2_X1 U108 ( .A(data_in[85]), .B(n827), .Z(n878) );
  XOR2_X1 U109 ( .A(data_in[69]), .B(data_in[93]), .Z(n827) );
  XOR2_X1 U110 ( .A(n879), .B(n880), .Z(data_out[76]) );
  XOR2_X1 U111 ( .A(n862), .B(n881), .Z(n880) );
  XOR2_X1 U112 ( .A(data_in[84]), .B(n830), .Z(n879) );
  XOR2_X1 U113 ( .A(data_in[68]), .B(data_in[92]), .Z(n830) );
  XOR2_X1 U114 ( .A(n882), .B(n883), .Z(data_out[75]) );
  XOR2_X1 U115 ( .A(n838), .B(n865), .Z(n883) );
  XOR2_X1 U116 ( .A(data_in[91]), .B(n884), .Z(n865) );
  XOR2_X1 U117 ( .A(data_in[87]), .B(data_in[82]), .Z(n884) );
  XOR2_X1 U118 ( .A(n885), .B(n886), .Z(data_out[74]) );
  XOR2_X1 U119 ( .A(data_in[66]), .B(n848), .Z(n886) );
  XOR2_X1 U120 ( .A(n887), .B(n888), .Z(data_out[73]) );
  XOR2_X1 U121 ( .A(n870), .B(n889), .Z(n888) );
  XOR2_X1 U122 ( .A(data_in[80]), .B(data_in[87]), .Z(n870) );
  XOR2_X1 U123 ( .A(data_in[81]), .B(n840), .Z(n887) );
  XOR2_X1 U124 ( .A(data_in[65]), .B(data_in[89]), .Z(n840) );
  XOR2_X1 U125 ( .A(n890), .B(n891), .Z(data_out[72]) );
  XOR2_X1 U126 ( .A(data_in[64]), .B(n892), .Z(n891) );
  XOR2_X1 U127 ( .A(data_in[87]), .B(data_in[79]), .Z(n890) );
  XOR2_X1 U128 ( .A(n893), .B(n894), .Z(data_out[71]) );
  XOR2_X1 U129 ( .A(data_in[70]), .B(n871), .Z(n894) );
  XOR2_X1 U130 ( .A(data_in[87]), .B(data_in[95]), .Z(n871) );
  XOR2_X1 U131 ( .A(data_in[79]), .B(data_in[78]), .Z(n893) );
  XOR2_X1 U132 ( .A(n895), .B(n896), .Z(data_out[70]) );
  XOR2_X1 U133 ( .A(data_in[69]), .B(n825), .Z(n896) );
  XOR2_X1 U134 ( .A(data_in[78]), .B(data_in[86]), .Z(n825) );
  XOR2_X1 U135 ( .A(data_in[94]), .B(data_in[77]), .Z(n895) );
  XOR2_X1 U136 ( .A(n897), .B(n898), .Z(data_out[6]) );
  XOR2_X1 U137 ( .A(data_in[13]), .B(n899), .Z(n898) );
  XOR2_X1 U138 ( .A(data_in[5]), .B(data_in[30]), .Z(n897) );
  XOR2_X1 U139 ( .A(n900), .B(n901), .Z(data_out[69]) );
  XOR2_X1 U140 ( .A(data_in[68]), .B(n828), .Z(n901) );
  XOR2_X1 U141 ( .A(data_in[77]), .B(data_in[85]), .Z(n828) );
  XOR2_X1 U142 ( .A(data_in[93]), .B(data_in[76]), .Z(n900) );
  XOR2_X1 U143 ( .A(n902), .B(n903), .Z(data_out[68]) );
  XOR2_X1 U144 ( .A(n834), .B(n881), .Z(n903) );
  XOR2_X1 U145 ( .A(data_in[75]), .B(data_in[79]), .Z(n881) );
  XOR2_X1 U146 ( .A(data_in[67]), .B(data_in[71]), .Z(n834) );
  XOR2_X1 U147 ( .A(data_in[92]), .B(n833), .Z(n902) );
  XOR2_X1 U148 ( .A(data_in[76]), .B(data_in[84]), .Z(n833) );
  XOR2_X1 U149 ( .A(n904), .B(n905), .Z(data_out[67]) );
  XOR2_X1 U150 ( .A(n839), .B(n882), .Z(n905) );
  XOR2_X1 U152 ( .A(data_in[71]), .B(data_in[66]), .Z(n906) );
  XOR2_X1 U153 ( .A(data_in[83]), .B(data_in[91]), .Z(n904) );
  XOR2_X1 U154 ( .A(n907), .B(n908), .Z(data_out[66]) );
  XOR2_X1 U155 ( .A(data_in[74]), .B(n885), .Z(n908) );
  XOR2_X1 U156 ( .A(data_in[90]), .B(data_in[82]), .Z(n885) );
  XOR2_X1 U157 ( .A(data_in[73]), .B(data_in[65]), .Z(n907) );
  XOR2_X1 U158 ( .A(n909), .B(n910), .Z(data_out[65]) );
  XOR2_X1 U159 ( .A(n849), .B(n889), .Z(n910) );
  XOR2_X1 U160 ( .A(data_in[72]), .B(data_in[79]), .Z(n889) );
  XOR2_X1 U161 ( .A(data_in[64]), .B(data_in[71]), .Z(n849) );
  XOR2_X1 U162 ( .A(data_in[89]), .B(n848), .Z(n909) );
  XOR2_X1 U163 ( .A(data_in[73]), .B(data_in[81]), .Z(n848) );
  XOR2_X1 U164 ( .A(n892), .B(n911), .Z(data_out[64]) );
  XOR2_X1 U165 ( .A(data_in[72]), .B(n822), .Z(n911) );
  XOR2_X1 U166 ( .A(data_in[71]), .B(data_in[79]), .Z(n822) );
  XOR2_X1 U167 ( .A(data_in[88]), .B(data_in[80]), .Z(n892) );
  XOR2_X1 U168 ( .A(n912), .B(n913), .Z(data_out[63]) );
  XOR2_X1 U169 ( .A(data_in[55]), .B(n914), .Z(n913) );
  XOR2_X1 U170 ( .A(n915), .B(n916), .Z(data_out[62]) );
  XOR2_X1 U171 ( .A(data_in[38]), .B(n917), .Z(n916) );
  XOR2_X1 U172 ( .A(n918), .B(n919), .Z(data_out[61]) );
  XOR2_X1 U173 ( .A(data_in[37]), .B(n920), .Z(n919) );
  XOR2_X1 U174 ( .A(n921), .B(n922), .Z(data_out[60]) );
  XOR2_X1 U175 ( .A(n923), .B(n924), .Z(n922) );
  XOR2_X1 U176 ( .A(data_in[36]), .B(n925), .Z(n921) );
  XOR2_X1 U177 ( .A(n926), .B(n927), .Z(data_out[5]) );
  XOR2_X1 U178 ( .A(data_in[12]), .B(n928), .Z(n927) );
  XOR2_X1 U179 ( .A(data_in[4]), .B(data_in[29]), .Z(n926) );
  XOR2_X1 U182 ( .A(n933), .B(n934), .Z(data_out[58]) );
  XOR2_X1 U183 ( .A(data_in[50]), .B(n935), .Z(n934) );
  XOR2_X1 U184 ( .A(n936), .B(n937), .Z(data_out[57]) );
  XOR2_X1 U185 ( .A(n938), .B(n939), .Z(n937) );
  XOR2_X1 U186 ( .A(data_in[33]), .B(n940), .Z(n936) );
  XOR2_X1 U187 ( .A(n941), .B(n942), .Z(data_out[56]) );
  XOR2_X1 U188 ( .A(data_in[48]), .B(n943), .Z(n942) );
  XOR2_X1 U189 ( .A(data_in[63]), .B(data_in[39]), .Z(n941) );
  XOR2_X1 U190 ( .A(n944), .B(n945), .Z(data_out[55]) );
  XOR2_X1 U191 ( .A(data_in[54]), .B(n912), .Z(n945) );
  XOR2_X1 U192 ( .A(data_in[63]), .B(data_in[62]), .Z(n944) );
  XOR2_X1 U193 ( .A(n946), .B(n947), .Z(data_out[54]) );
  XOR2_X1 U194 ( .A(data_in[46]), .B(n914), .Z(n947) );
  XOR2_X1 U195 ( .A(data_in[61]), .B(data_in[53]), .Z(n946) );
  XOR2_X1 U196 ( .A(n948), .B(n949), .Z(data_out[53]) );
  XOR2_X1 U197 ( .A(data_in[45]), .B(n917), .Z(n949) );
  XOR2_X1 U198 ( .A(data_in[60]), .B(data_in[52]), .Z(n948) );
  XOR2_X1 U199 ( .A(n950), .B(n951), .Z(data_out[52]) );
  XOR2_X1 U200 ( .A(n925), .B(n952), .Z(n951) );
  XOR2_X1 U201 ( .A(data_in[59]), .B(data_in[63]), .Z(n925) );
  XOR2_X1 U202 ( .A(data_in[44]), .B(n920), .Z(n950) );
  XOR2_X1 U203 ( .A(n953), .B(n954), .Z(data_out[51]) );
  XOR2_X1 U204 ( .A(data_in[58]), .B(data_in[63]), .Z(n930) );
  XOR2_X1 U205 ( .A(n956), .B(n957), .Z(data_out[50]) );
  XOR2_X1 U206 ( .A(data_in[58]), .B(n935), .Z(n957) );
  XOR2_X1 U207 ( .A(data_in[42]), .B(data_in[34]), .Z(n935) );
  XOR2_X1 U208 ( .A(data_in[57]), .B(data_in[49]), .Z(n956) );
  XOR2_X1 U209 ( .A(n958), .B(n959), .Z(data_out[4]) );
  XOR2_X1 U210 ( .A(n960), .B(n961), .Z(n959) );
  XOR2_X1 U211 ( .A(data_in[28]), .B(n962), .Z(n958) );
  XOR2_X1 U212 ( .A(n963), .B(n964), .Z(data_out[49]) );
  XOR2_X1 U213 ( .A(n940), .B(n965), .Z(n964) );
  XOR2_X1 U214 ( .A(data_in[56]), .B(data_in[63]), .Z(n940) );
  XOR2_X1 U215 ( .A(data_in[41]), .B(n933), .Z(n963) );
  XOR2_X1 U216 ( .A(n966), .B(n967), .Z(data_out[48]) );
  XOR2_X1 U217 ( .A(data_in[56]), .B(n943), .Z(n967) );
  XOR2_X1 U218 ( .A(data_in[40]), .B(data_in[32]), .Z(n943) );
  XOR2_X1 U219 ( .A(n966), .B(n968), .Z(data_out[47]) );
  XOR2_X1 U220 ( .A(data_in[39]), .B(n915), .Z(n968) );
  XOR2_X1 U221 ( .A(n918), .B(n969), .Z(data_out[46]) );
  XOR2_X1 U222 ( .A(data_in[54]), .B(n914), .Z(n969) );
  XOR2_X1 U223 ( .A(data_in[38]), .B(data_in[62]), .Z(n914) );
  XOR2_X1 U224 ( .A(n923), .B(n970), .Z(data_out[45]) );
  XOR2_X1 U225 ( .A(data_in[53]), .B(n917), .Z(n970) );
  XOR2_X1 U226 ( .A(data_in[37]), .B(data_in[61]), .Z(n917) );
  XOR2_X1 U227 ( .A(n971), .B(n972), .Z(data_out[44]) );
  XOR2_X1 U228 ( .A(n952), .B(n973), .Z(n972) );
  XOR2_X1 U229 ( .A(data_in[52]), .B(n920), .Z(n971) );
  XOR2_X1 U230 ( .A(data_in[36]), .B(data_in[60]), .Z(n920) );
  XOR2_X1 U231 ( .A(n974), .B(n975), .Z(data_out[43]) );
  XOR2_X1 U232 ( .A(n931), .B(n955), .Z(n975) );
  XOR2_X1 U233 ( .A(data_in[59]), .B(n976), .Z(n955) );
  XOR2_X1 U234 ( .A(data_in[55]), .B(data_in[50]), .Z(n976) );
  XOR2_X1 U235 ( .A(n977), .B(n978), .Z(data_out[42]) );
  XOR2_X1 U236 ( .A(data_in[34]), .B(n938), .Z(n978) );
  XOR2_X1 U237 ( .A(n979), .B(n980), .Z(data_out[41]) );
  XOR2_X1 U238 ( .A(n965), .B(n981), .Z(n980) );
  XOR2_X1 U239 ( .A(data_in[48]), .B(data_in[55]), .Z(n965) );
  XOR2_X1 U240 ( .A(data_in[49]), .B(n933), .Z(n979) );
  XOR2_X1 U241 ( .A(data_in[33]), .B(data_in[57]), .Z(n933) );
  XOR2_X1 U242 ( .A(n982), .B(n983), .Z(data_out[40]) );
  XOR2_X1 U243 ( .A(data_in[32]), .B(n984), .Z(n983) );
  XOR2_X1 U244 ( .A(data_in[55]), .B(data_in[47]), .Z(n982) );
  XOR2_X1 U245 ( .A(n985), .B(n986), .Z(data_out[3]) );
  XOR2_X1 U246 ( .A(data_in[19]), .B(data_in[27]), .Z(n985) );
  XOR2_X1 U247 ( .A(n989), .B(n990), .Z(data_out[39]) );
  XOR2_X1 U248 ( .A(data_in[38]), .B(n966), .Z(n990) );
  XOR2_X1 U249 ( .A(data_in[55]), .B(data_in[63]), .Z(n966) );
  XOR2_X1 U250 ( .A(data_in[47]), .B(data_in[46]), .Z(n989) );
  XOR2_X1 U251 ( .A(n991), .B(n992), .Z(data_out[38]) );
  XOR2_X1 U252 ( .A(data_in[37]), .B(n915), .Z(n992) );
  XOR2_X1 U253 ( .A(data_in[46]), .B(data_in[54]), .Z(n915) );
  XOR2_X1 U254 ( .A(data_in[62]), .B(data_in[45]), .Z(n991) );
  XOR2_X1 U255 ( .A(n993), .B(n994), .Z(data_out[37]) );
  XOR2_X1 U256 ( .A(data_in[36]), .B(n918), .Z(n994) );
  XOR2_X1 U257 ( .A(data_in[45]), .B(data_in[53]), .Z(n918) );
  XOR2_X1 U258 ( .A(data_in[61]), .B(data_in[44]), .Z(n993) );
  XOR2_X1 U259 ( .A(n995), .B(n996), .Z(data_out[36]) );
  XOR2_X1 U260 ( .A(n924), .B(n973), .Z(n996) );
  XOR2_X1 U261 ( .A(data_in[43]), .B(data_in[47]), .Z(n973) );
  XOR2_X1 U262 ( .A(data_in[35]), .B(data_in[39]), .Z(n924) );
  XOR2_X1 U263 ( .A(data_in[60]), .B(n923), .Z(n995) );
  XOR2_X1 U264 ( .A(data_in[44]), .B(data_in[52]), .Z(n923) );
  XOR2_X1 U265 ( .A(n997), .B(n998), .Z(data_out[35]) );
  XOR2_X1 U266 ( .A(n932), .B(n974), .Z(n998) );
  XOR2_X1 U268 ( .A(data_in[39]), .B(data_in[34]), .Z(n999) );
  XOR2_X1 U269 ( .A(data_in[51]), .B(data_in[59]), .Z(n997) );
  XOR2_X1 U270 ( .A(n1000), .B(n1001), .Z(data_out[34]) );
  XOR2_X1 U271 ( .A(data_in[42]), .B(n977), .Z(n1001) );
  XOR2_X1 U272 ( .A(data_in[58]), .B(data_in[50]), .Z(n977) );
  XOR2_X1 U273 ( .A(data_in[41]), .B(data_in[33]), .Z(n1000) );
  XOR2_X1 U274 ( .A(n1002), .B(n1003), .Z(data_out[33]) );
  XOR2_X1 U275 ( .A(n939), .B(n981), .Z(n1003) );
  XOR2_X1 U276 ( .A(data_in[40]), .B(data_in[47]), .Z(n981) );
  XOR2_X1 U277 ( .A(data_in[32]), .B(data_in[39]), .Z(n939) );
  XOR2_X1 U278 ( .A(data_in[57]), .B(n938), .Z(n1002) );
  XOR2_X1 U279 ( .A(data_in[41]), .B(data_in[49]), .Z(n938) );
  XOR2_X1 U280 ( .A(n984), .B(n1004), .Z(data_out[32]) );
  XOR2_X1 U281 ( .A(data_in[40]), .B(n912), .Z(n1004) );
  XOR2_X1 U282 ( .A(data_in[39]), .B(data_in[47]), .Z(n912) );
  XOR2_X1 U283 ( .A(data_in[56]), .B(data_in[48]), .Z(n984) );
  XOR2_X1 U284 ( .A(n1005), .B(n1006), .Z(data_out[31]) );
  XOR2_X1 U285 ( .A(data_in[23]), .B(n1007), .Z(n1006) );
  XOR2_X1 U286 ( .A(n1008), .B(n1009), .Z(data_out[30]) );
  XOR2_X1 U287 ( .A(data_in[6]), .B(n899), .Z(n1009) );
  XOR2_X1 U288 ( .A(n1010), .B(n1011), .Z(data_out[2]) );
  XOR2_X1 U289 ( .A(data_in[10]), .B(n1012), .Z(n1011) );
  XOR2_X1 U290 ( .A(data_in[9]), .B(data_in[1]), .Z(n1010) );
  XOR2_X1 U291 ( .A(n1013), .B(n1014), .Z(data_out[29]) );
  XOR2_X1 U292 ( .A(data_in[5]), .B(n928), .Z(n1014) );
  XOR2_X1 U293 ( .A(n1015), .B(n1016), .Z(data_out[28]) );
  XOR2_X1 U294 ( .A(n960), .B(n1017), .Z(n1016) );
  XOR2_X1 U295 ( .A(data_in[3]), .B(data_in[7]), .Z(n960) );
  XOR2_X1 U296 ( .A(data_in[4]), .B(n962), .Z(n1015) );
  XOR2_X1 U298 ( .A(data_in[7]), .B(data_in[2]), .Z(n1020) );
  XOR2_X1 U299 ( .A(n1022), .B(n1023), .Z(data_out[26]) );
  XOR2_X1 U300 ( .A(data_in[18]), .B(n806), .Z(n1023) );
  XOR2_X1 U301 ( .A(n1024), .B(n1025), .Z(data_out[25]) );
  XOR2_X1 U302 ( .A(data_in[1]), .B(n1026), .Z(n1024) );
  XOR2_X1 U303 ( .A(n1027), .B(n1028), .Z(data_out[24]) );
  XOR2_X1 U304 ( .A(data_in[16]), .B(n1029), .Z(n1028) );
  XOR2_X1 U305 ( .A(data_in[7]), .B(data_in[31]), .Z(n1027) );
  XOR2_X1 U306 ( .A(n1030), .B(n1031), .Z(data_out[23]) );
  XOR2_X1 U307 ( .A(data_in[22]), .B(n1005), .Z(n1031) );
  XOR2_X1 U308 ( .A(data_in[31]), .B(data_in[30]), .Z(n1030) );
  XOR2_X1 U309 ( .A(n1032), .B(n1033), .Z(data_out[22]) );
  XOR2_X1 U310 ( .A(data_in[14]), .B(n1007), .Z(n1033) );
  XOR2_X1 U311 ( .A(data_in[29]), .B(data_in[21]), .Z(n1032) );
  XOR2_X1 U312 ( .A(n1034), .B(n1035), .Z(data_out[21]) );
  XOR2_X1 U313 ( .A(data_in[13]), .B(n1008), .Z(n1035) );
  XOR2_X1 U314 ( .A(data_in[28]), .B(data_in[20]), .Z(n1034) );
  XOR2_X1 U315 ( .A(n1036), .B(n1037), .Z(data_out[20]) );
  XOR2_X1 U316 ( .A(n1017), .B(n1038), .Z(n1037) );
  XOR2_X1 U317 ( .A(data_in[27]), .B(data_in[31]), .Z(n1017) );
  XOR2_X1 U318 ( .A(data_in[12]), .B(n1013), .Z(n1036) );
  XOR2_X1 U319 ( .A(n1039), .B(n1025), .Z(data_out[1]) );
  XOR2_X1 U320 ( .A(n1040), .B(n1041), .Z(n1025) );
  XOR2_X1 U321 ( .A(data_in[0]), .B(data_in[7]), .Z(n1041) );
  XOR2_X1 U322 ( .A(data_in[25]), .B(n805), .Z(n1039) );
  XOR2_X1 U323 ( .A(data_in[8]), .B(data_in[15]), .Z(n805) );
  XOR2_X1 U324 ( .A(n1042), .B(n1043), .Z(data_out[19]) );
  XOR2_X1 U325 ( .A(n1021), .B(n1044), .Z(n1043) );
  XOR2_X1 U327 ( .A(n1045), .B(n1046), .Z(data_out[18]) );
  XOR2_X1 U328 ( .A(data_in[26]), .B(n1022), .Z(n1046) );
  XOR2_X1 U329 ( .A(data_in[10]), .B(data_in[2]), .Z(n1022) );
  XOR2_X1 U330 ( .A(data_in[25]), .B(data_in[17]), .Z(n1045) );
  XOR2_X1 U331 ( .A(n1047), .B(n1048), .Z(data_out[17]) );
  XOR2_X1 U332 ( .A(n804), .B(n1026), .Z(n1048) );
  XOR2_X1 U333 ( .A(data_in[24]), .B(data_in[31]), .Z(n1026) );
  XOR2_X1 U334 ( .A(data_in[16]), .B(data_in[23]), .Z(n804) );
  XOR2_X1 U335 ( .A(data_in[9]), .B(n806), .Z(n1047) );
  XOR2_X1 U336 ( .A(data_in[1]), .B(data_in[25]), .Z(n806) );
  XOR2_X1 U337 ( .A(n1029), .B(n1049), .Z(data_out[16]) );
  XOR2_X1 U338 ( .A(data_in[24]), .B(n875), .Z(n1049) );
  XOR2_X1 U339 ( .A(data_in[8]), .B(data_in[0]), .Z(n1029) );
  XOR2_X1 U340 ( .A(n899), .B(n1050), .Z(data_out[15]) );
  XOR2_X1 U341 ( .A(data_in[7]), .B(n875), .Z(n1050) );
  XOR2_X1 U342 ( .A(data_in[23]), .B(data_in[31]), .Z(n875) );
  XOR2_X1 U343 ( .A(data_in[14]), .B(data_in[22]), .Z(n899) );
  XOR2_X1 U344 ( .A(n1007), .B(n1051), .Z(data_out[14]) );
  XOR2_X1 U345 ( .A(data_in[22]), .B(n928), .Z(n1051) );
  XOR2_X1 U346 ( .A(data_in[13]), .B(data_in[21]), .Z(n928) );
  XOR2_X1 U347 ( .A(data_in[30]), .B(data_in[6]), .Z(n1007) );
  XOR2_X1 U348 ( .A(n1008), .B(n1052), .Z(data_out[13]) );
  XOR2_X1 U349 ( .A(data_in[21]), .B(n962), .Z(n1052) );
  XOR2_X1 U350 ( .A(data_in[12]), .B(data_in[20]), .Z(n962) );
  XOR2_X1 U351 ( .A(data_in[29]), .B(data_in[5]), .Z(n1008) );
  XOR2_X1 U352 ( .A(n1053), .B(n1054), .Z(data_out[12]) );
  XOR2_X1 U353 ( .A(n1013), .B(n1038), .Z(n1054) );
  XOR2_X1 U354 ( .A(data_in[19]), .B(data_in[23]), .Z(n1038) );
  XOR2_X1 U355 ( .A(data_in[28]), .B(data_in[4]), .Z(n1013) );
  XOR2_X1 U356 ( .A(data_in[20]), .B(n961), .Z(n1053) );
  XOR2_X1 U357 ( .A(data_in[11]), .B(data_in[15]), .Z(n961) );
  XOR2_X1 U358 ( .A(n1055), .B(n1056), .Z(data_out[127]) );
  XOR2_X1 U359 ( .A(data_in[119]), .B(n819), .Z(n1056) );
  XOR2_X1 U360 ( .A(n1057), .B(n1058), .Z(data_out[126]) );
  XOR2_X1 U361 ( .A(data_in[102]), .B(n1059), .Z(n1058) );
  XOR2_X1 U362 ( .A(n1060), .B(n1061), .Z(data_out[125]) );
  XOR2_X1 U363 ( .A(data_in[101]), .B(n1062), .Z(n1061) );
  XOR2_X1 U364 ( .A(n1063), .B(n1064), .Z(data_out[124]) );
  XOR2_X1 U365 ( .A(n1065), .B(n1066), .Z(n1064) );
  XOR2_X1 U366 ( .A(data_in[100]), .B(n1067), .Z(n1063) );
  XOR2_X1 U368 ( .A(data_in[103]), .B(data_in[98]), .Z(n1070) );
  XOR2_X1 U369 ( .A(n1072), .B(n1073), .Z(data_out[122]) );
  XOR2_X1 U370 ( .A(data_in[114]), .B(n1074), .Z(n1073) );
  XOR2_X1 U371 ( .A(n1075), .B(n1076), .Z(data_out[121]) );
  XOR2_X1 U372 ( .A(n817), .B(n1077), .Z(n1076) );
  XOR2_X1 U373 ( .A(data_in[97]), .B(n818), .Z(n1075) );
  XOR2_X1 U374 ( .A(n1078), .B(n1079), .Z(data_out[120]) );
  XOR2_X1 U375 ( .A(data_in[112]), .B(n1080), .Z(n1079) );
  XOR2_X1 U376 ( .A(data_in[127]), .B(data_in[103]), .Z(n1078) );
  XOR2_X1 U377 ( .A(n1044), .B(n1081), .Z(data_out[11]) );
  XOR2_X1 U378 ( .A(n988), .B(n1019), .Z(n1081) );
  XOR2_X1 U379 ( .A(data_in[10]), .B(data_in[15]), .Z(n988) );
  XOR2_X1 U380 ( .A(data_in[27]), .B(n1082), .Z(n1044) );
  XOR2_X1 U381 ( .A(data_in[23]), .B(data_in[18]), .Z(n1082) );
  XOR2_X1 U382 ( .A(n1083), .B(n1084), .Z(data_out[119]) );
  XOR2_X1 U383 ( .A(data_in[118]), .B(n819), .Z(n1084) );
  XOR2_X1 U384 ( .A(data_in[103]), .B(data_in[111]), .Z(n819) );
  XOR2_X1 U385 ( .A(data_in[127]), .B(data_in[126]), .Z(n1083) );
  XOR2_X1 U386 ( .A(n1085), .B(n1086), .Z(data_out[118]) );
  XOR2_X1 U387 ( .A(data_in[110]), .B(n1055), .Z(n1086) );
  XOR2_X1 U388 ( .A(data_in[125]), .B(data_in[117]), .Z(n1085) );
  XOR2_X1 U389 ( .A(n1087), .B(n1088), .Z(data_out[117]) );
  XOR2_X1 U390 ( .A(data_in[109]), .B(n1059), .Z(n1088) );
  XOR2_X1 U391 ( .A(data_in[124]), .B(data_in[116]), .Z(n1087) );
  XOR2_X1 U392 ( .A(n1089), .B(n1090), .Z(data_out[116]) );
  XOR2_X1 U393 ( .A(n1067), .B(n1091), .Z(n1090) );
  XOR2_X1 U394 ( .A(data_in[123]), .B(data_in[127]), .Z(n1067) );
  XOR2_X1 U395 ( .A(data_in[108]), .B(n1062), .Z(n1089) );
  XOR2_X1 U396 ( .A(n1092), .B(n1093), .Z(data_out[115]) );
  XOR2_X1 U397 ( .A(n1071), .B(n1094), .Z(n1093) );
  XOR2_X1 U399 ( .A(n1095), .B(n1096), .Z(data_out[114]) );
  XOR2_X1 U400 ( .A(data_in[122]), .B(n1074), .Z(n1096) );
  XOR2_X1 U401 ( .A(data_in[106]), .B(data_in[98]), .Z(n1074) );
  XOR2_X1 U402 ( .A(data_in[121]), .B(data_in[113]), .Z(n1095) );
  XOR2_X1 U403 ( .A(n1097), .B(n1098), .Z(data_out[113]) );
  XOR2_X1 U404 ( .A(n1077), .B(n1099), .Z(n1098) );
  XOR2_X1 U405 ( .A(data_in[120]), .B(data_in[127]), .Z(n1077) );
  XOR2_X1 U406 ( .A(data_in[105]), .B(n1072), .Z(n1097) );
  XOR2_X1 U407 ( .A(n1100), .B(n1101), .Z(data_out[112]) );
  XOR2_X1 U408 ( .A(data_in[120]), .B(n1080), .Z(n1101) );
  XOR2_X1 U409 ( .A(data_in[104]), .B(data_in[96]), .Z(n1080) );
  XOR2_X1 U410 ( .A(n1100), .B(n1102), .Z(data_out[111]) );
  XOR2_X1 U411 ( .A(data_in[103]), .B(n1057), .Z(n1102) );
  XOR2_X1 U412 ( .A(n1060), .B(n1103), .Z(data_out[110]) );
  XOR2_X1 U413 ( .A(data_in[118]), .B(n1055), .Z(n1103) );
  XOR2_X1 U414 ( .A(data_in[102]), .B(data_in[126]), .Z(n1055) );
  XOR2_X1 U415 ( .A(n1040), .B(n1104), .Z(data_out[10]) );
  XOR2_X1 U416 ( .A(data_in[2]), .B(n1012), .Z(n1104) );
  XOR2_X1 U417 ( .A(data_in[26]), .B(data_in[18]), .Z(n1012) );
  XOR2_X1 U418 ( .A(data_in[17]), .B(data_in[9]), .Z(n1040) );
  XOR2_X1 U419 ( .A(n1065), .B(n1105), .Z(data_out[109]) );
  XOR2_X1 U420 ( .A(data_in[117]), .B(n1059), .Z(n1105) );
  XOR2_X1 U421 ( .A(data_in[101]), .B(data_in[125]), .Z(n1059) );
  XOR2_X1 U422 ( .A(n1106), .B(n1107), .Z(data_out[108]) );
  XOR2_X1 U423 ( .A(n1091), .B(n1108), .Z(n1107) );
  XOR2_X1 U424 ( .A(data_in[115]), .B(data_in[119]), .Z(n1091) );
  XOR2_X1 U425 ( .A(data_in[116]), .B(n1062), .Z(n1106) );
  XOR2_X1 U426 ( .A(data_in[100]), .B(data_in[124]), .Z(n1062) );
  XOR2_X1 U427 ( .A(n1094), .B(n1109), .Z(data_out[107]) );
  XOR2_X1 U428 ( .A(n810), .B(n1069), .Z(n1109) );
  XOR2_X1 U429 ( .A(data_in[106]), .B(data_in[111]), .Z(n810) );
  XOR2_X1 U430 ( .A(data_in[123]), .B(n1110), .Z(n1094) );
  XOR2_X1 U431 ( .A(data_in[119]), .B(data_in[114]), .Z(n1110) );
  XOR2_X1 U432 ( .A(n818), .B(n1111), .Z(data_out[106]) );
  XOR2_X1 U433 ( .A(data_in[98]), .B(n813), .Z(n1111) );
  XOR2_X1 U434 ( .A(data_in[122]), .B(data_in[114]), .Z(n813) );
  XOR2_X1 U435 ( .A(data_in[105]), .B(data_in[113]), .Z(n818) );
  XOR2_X1 U436 ( .A(n1112), .B(n1113), .Z(data_out[105]) );
  XOR2_X1 U437 ( .A(n1072), .B(n1099), .Z(n1113) );
  XOR2_X1 U438 ( .A(data_in[112]), .B(data_in[119]), .Z(n1099) );
  XOR2_X1 U439 ( .A(data_in[121]), .B(data_in[97]), .Z(n1072) );
  XOR2_X1 U440 ( .A(data_in[113]), .B(n816), .Z(n1112) );
  XOR2_X1 U441 ( .A(data_in[104]), .B(data_in[111]), .Z(n816) );
  XOR2_X1 U442 ( .A(n1114), .B(n1115), .Z(data_out[104]) );
  XOR2_X1 U443 ( .A(data_in[96]), .B(n821), .Z(n1115) );
  XOR2_X1 U444 ( .A(data_in[120]), .B(data_in[112]), .Z(n821) );
  XOR2_X1 U445 ( .A(data_in[119]), .B(data_in[111]), .Z(n1114) );
  XOR2_X1 U446 ( .A(n1116), .B(n1117), .Z(data_out[103]) );
  XOR2_X1 U447 ( .A(data_in[102]), .B(n1100), .Z(n1117) );
  XOR2_X1 U448 ( .A(data_in[119]), .B(data_in[127]), .Z(n1100) );
  XOR2_X1 U449 ( .A(data_in[111]), .B(data_in[110]), .Z(n1116) );
  XOR2_X1 U450 ( .A(n1118), .B(n1119), .Z(data_out[102]) );
  XOR2_X1 U451 ( .A(data_in[101]), .B(n1057), .Z(n1119) );
  XOR2_X1 U452 ( .A(data_in[110]), .B(data_in[118]), .Z(n1057) );
  XOR2_X1 U453 ( .A(data_in[126]), .B(data_in[109]), .Z(n1118) );
  XOR2_X1 U454 ( .A(n1120), .B(n1121), .Z(data_out[101]) );
  XOR2_X1 U455 ( .A(data_in[100]), .B(n1060), .Z(n1121) );
  XOR2_X1 U456 ( .A(data_in[109]), .B(data_in[117]), .Z(n1060) );
  XOR2_X1 U457 ( .A(data_in[125]), .B(data_in[108]), .Z(n1120) );
  XOR2_X1 U458 ( .A(n1122), .B(n1123), .Z(data_out[100]) );
  XOR2_X1 U459 ( .A(n1066), .B(n1108), .Z(n1123) );
  XOR2_X1 U460 ( .A(data_in[107]), .B(data_in[111]), .Z(n1108) );
  XOR2_X1 U461 ( .A(data_in[124]), .B(n1065), .Z(n1122) );
  XOR2_X1 U462 ( .A(data_in[108]), .B(data_in[116]), .Z(n1065) );
  XOR2_X1 U463 ( .A(n1005), .B(n1124), .Z(data_out[0]) );
  XOR2_X1 U464 ( .A(data_in[8]), .B(n845), .Z(n1124) );
  XOR2_X1 U465 ( .A(data_in[24]), .B(data_in[16]), .Z(n845) );
  XOR2_X1 U466 ( .A(data_in[15]), .B(data_in[7]), .Z(n1005) );
  INV_X1 U467 ( .A(n931), .ZN(n796) );
  INV_X1 U468 ( .A(n838), .ZN(n792) );
  XOR2_X1 U469 ( .A(n1021), .B(n1125), .Z(data_out[27]) );
  XOR2_X1 U470 ( .A(n987), .B(n1019), .Z(n1125) );
  XOR2_X1 U471 ( .A(n932), .B(n1126), .Z(data_out[59]) );
  XNOR2_X1 U472 ( .A(n796), .B(n930), .ZN(n1126) );
  XOR2_X1 U473 ( .A(n839), .B(n1127), .Z(data_out[91]) );
  XNOR2_X1 U474 ( .A(n792), .B(n837), .ZN(n1127) );
  XOR2_X1 U475 ( .A(n1071), .B(n1128), .Z(data_out[123]) );
  XOR2_X1 U476 ( .A(n809), .B(n1069), .Z(n1128) );
  XNOR2_X1 U477 ( .A(data_in[26]), .B(data_in[31]), .ZN(n1021) );
  XNOR2_X1 U478 ( .A(data_in[122]), .B(data_in[127]), .ZN(n1071) );
  XNOR2_X1 U479 ( .A(data_in[42]), .B(data_in[47]), .ZN(n974) );
  XNOR2_X1 U480 ( .A(data_in[74]), .B(data_in[79]), .ZN(n882) );
  XNOR2_X1 U481 ( .A(data_in[11]), .B(data_in[3]), .ZN(n1042) );
  XNOR2_X1 U482 ( .A(data_in[43]), .B(data_in[35]), .ZN(n953) );
  XNOR2_X1 U483 ( .A(n930), .B(n955), .ZN(n954) );
  XNOR2_X1 U484 ( .A(data_in[75]), .B(data_in[67]), .ZN(n863) );
  XNOR2_X1 U485 ( .A(n837), .B(n865), .ZN(n864) );
  XNOR2_X1 U486 ( .A(data_in[107]), .B(data_in[99]), .ZN(n1092) );
  XNOR2_X1 U487 ( .A(n987), .B(n988), .ZN(n986) );
  XNOR2_X1 U488 ( .A(data_in[11]), .B(n1020), .ZN(n987) );
  XNOR2_X1 U489 ( .A(data_in[107]), .B(n1070), .ZN(n809) );
  XOR2_X1 U490 ( .A(data_in[115]), .B(data_in[99]), .Z(n1069) );
  XOR2_X1 U491 ( .A(data_in[19]), .B(data_in[3]), .Z(n1019) );
  XNOR2_X1 U492 ( .A(data_in[43]), .B(n999), .ZN(n932) );
  XNOR2_X1 U493 ( .A(data_in[75]), .B(n906), .ZN(n839) );
  XNOR2_X1 U494 ( .A(data_in[51]), .B(data_in[35]), .ZN(n931) );
  XNOR2_X1 U495 ( .A(data_in[83]), .B(data_in[67]), .ZN(n838) );
  XNOR2_X1 U496 ( .A(data_in[96]), .B(n790), .ZN(n817) );
  XNOR2_X1 U497 ( .A(data_in[99]), .B(n790), .ZN(n1066) );
  XOR2_X1 U498 ( .A(data_in[51]), .B(data_in[55]), .Z(n952) );
  XOR2_X1 U499 ( .A(data_in[83]), .B(data_in[87]), .Z(n862) );
  XNOR2_X1 U500 ( .A(n809), .B(n810), .ZN(n808) );
  INV_X1 U501 ( .A(data_in[103]), .ZN(n790) );
endmodule

